////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
/// TSMC Library/IP Product
/// Filename: tcbn65lpbwp12tlvt.v
/// Technology: CLN65LP
/// Product Type: Standard Cell
/// Product Name: tcbn65lpbwp12tlvt
/// Version: 140c
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////
///  STATEMENT OF USE
///
///  This information contains confidential and proprietary information of TSMC.
///  No part of this information may be reproduced, transmitted, transcribed,
///  stored in a retrieval system, or translated into any human or computer
///  language, in any form or by any means, electronic, mechanical, magnetic,
///  optical, chemical, manual, or otherwise, without the prior written permission
///  of TSMC.  This information was prepared for informational purpose and is for
///  use by TSMC's customers only.  TSMC reserves the right to make changes in the
///  information at any time and without notice.
///
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
`timescale 1ns/10ps

`celldefine
module AN2D0BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN2D1BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN2D2BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN2D4BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN2D8BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN2XD1BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN3D0BWP12TLVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    and		(Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN3D1BWP12TLVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    and		(Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN3D2BWP12TLVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    and		(Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN3D4BWP12TLVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    and		(Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN3D8BWP12TLVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    and		(Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN3XD1BWP12TLVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    and		(Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN4D0BWP12TLVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    and		(Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN4D1BWP12TLVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    and		(Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN4D2BWP12TLVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    and		(Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN4D4BWP12TLVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    and		(Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN4D8BWP12TLVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    and		(Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN4XD1BWP12TLVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    and		(Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ANTENNABWP12TLVT (I);
  input I;
  buf (I_buf, I);

endmodule
`endcelldefine

`celldefine
module AO211D0BWP12TLVT (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    and		(A, A1, A2);
    or		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B => Z) = (0, 0);
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO211D1BWP12TLVT (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    and		(A, A1, A2);
    or		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B => Z) = (0, 0);
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO211D2BWP12TLVT (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    and		(A, A1, A2);
    or		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B => Z) = (0, 0);
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO211D4BWP12TLVT (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    and		(A, A1, A2);
    or		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B => Z) = (0, 0);
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO21D0BWP12TLVT (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    and		(A, A1, A2);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO21D1BWP12TLVT (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    and		(A, A1, A2);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO21D2BWP12TLVT (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    and		(A, A1, A2);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO21D4BWP12TLVT (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    and		(A, A1, A2);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO221D0BWP12TLVT (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    and		(A, A1, A2);
    and     (B, B1, B2);
    or		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO221D1BWP12TLVT (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    and		(A, A1, A2);
    and     (B, B1, B2);
    or		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO221D2BWP12TLVT (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    and		(A, A1, A2);
    and     (B, B1, B2);
    or		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO221D4BWP12TLVT (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    and		(A, A1, A2);
    and     (B, B1, B2);
    or		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO222D0BWP12TLVT (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    and		(A, A1, A2);
    and     (B, B1, B2);
    and     (C, C1, C2);
    or		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (C1 => Z) = (0, 0);
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO222D1BWP12TLVT (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    and		(A, A1, A2);
    and     (B, B1, B2);
    and     (C, C1, C2);
    or		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (C1 => Z) = (0, 0);
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO222D2BWP12TLVT (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    and		(A, A1, A2);
    and     (B, B1, B2);
    and     (C, C1, C2);
    or		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (C1 => Z) = (0, 0);
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO222D4BWP12TLVT (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    and		(A, A1, A2);
    and     (B, B1, B2);
    and     (C, C1, C2);
    or		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (C1 => Z) = (0, 0);
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO22D0BWP12TLVT (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    and		(A, A1, A2);
    and     (B, B1, B2);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO22D1BWP12TLVT (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    and		(A, A1, A2);
    and     (B, B1, B2);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO22D2BWP12TLVT (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    and		(A, A1, A2);
    and     (B, B1, B2);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO22D4BWP12TLVT (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    and		(A, A1, A2);
    and     (B, B1, B2);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO31D0BWP12TLVT (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    and		(A, A1, A2, A3);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO31D1BWP12TLVT (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    and		(A, A1, A2, A3);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO31D2BWP12TLVT (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    and		(A, A1, A2, A3);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO31D4BWP12TLVT (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    and		(A, A1, A2, A3);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO32D0BWP12TLVT (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    and		(A, A1, A2, A3);
    and		(B, B1, B2);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO32D1BWP12TLVT (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    and		(A, A1, A2, A3);
    and		(B, B1, B2);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO32D2BWP12TLVT (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    and		(A, A1, A2, A3);
    and		(B, B1, B2);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO32D4BWP12TLVT (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    and		(A, A1, A2, A3);
    and		(B, B1, B2);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO33D0BWP12TLVT (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    and		(A, A1, A2, A3);
    and		(B, B1, B2, B3);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO33D1BWP12TLVT (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    and		(A, A1, A2, A3);
    and		(B, B1, B2, B3);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO33D2BWP12TLVT (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    and		(A, A1, A2, A3);
    and		(B, B1, B2, B3);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO33D4BWP12TLVT (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    and		(A, A1, A2, A3);
    and		(B, B1, B2, B3);
    or		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211D0BWP12TLVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and		(A, A1, A2);
    nor		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211D1BWP12TLVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and		(A, A1, A2);
    nor		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211D2BWP12TLVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and		(A, A1, A2);
    nor		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211D4BWP12TLVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and		(A, A1, A2);
    nor		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211XD0BWP12TLVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and		(A, A1, A2);
    nor		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211XD1BWP12TLVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and		(A, A1, A2);
    nor		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211XD2BWP12TLVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and		(A, A1, A2);
    nor		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211XD4BWP12TLVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and		(A, A1, A2);
    nor		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI21D0BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and		(A, A1, A2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI21D1BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and		(A, A1, A2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI21D2BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and		(A, A1, A2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI21D4BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and		(A, A1, A2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI221D0BWP12TLVT (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    and		(A, A1, A2);
    and		(B, B1, B2);
    nor		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI221D1BWP12TLVT (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    and		(A, A1, A2);
    and		(B, B1, B2);
    nor		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI221D2BWP12TLVT (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    and		(A, A1, A2);
    and		(B, B1, B2);
    nor		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI221D4BWP12TLVT (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    and		(A, A1, A2);
    and		(B, B1, B2);
    nor		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI221XD4BWP12TLVT (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    and		(A, A1, A2);
    and		(B, B1, B2);
    nor		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI222D0BWP12TLVT (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    and		(A, A1, A2);
    and		(B, B1, B2);
    and		(C, C1, C2);
    nor		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C1 => ZN) = (0, 0);
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI222D1BWP12TLVT (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    and		(A, A1, A2);
    and		(B, B1, B2);
    and		(C, C1, C2);
    nor		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C1 => ZN) = (0, 0);
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI222D2BWP12TLVT (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    and		(A, A1, A2);
    and		(B, B1, B2);
    and		(C, C1, C2);
    nor		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C1 => ZN) = (0, 0);
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI222D4BWP12TLVT (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    and		(A, A1, A2);
    and		(B, B1, B2);
    and		(C, C1, C2);
    nor		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C1 => ZN) = (0, 0);
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI222XD4BWP12TLVT (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    and		(A, A1, A2);
    and		(B, B1, B2);
    and		(C, C1, C2);
    nor		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C1 => ZN) = (0, 0);
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI22D0BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and		(A, A1, A2);
    and		(B, B1, B2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI22D1BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and		(A, A1, A2);
    and		(B, B1, B2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI22D2BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and		(A, A1, A2);
    and		(B, B1, B2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI22D4BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and		(A, A1, A2);
    and		(B, B1, B2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI31D0BWP12TLVT (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    and		(A, A1, A2, A3);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI31D1BWP12TLVT (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    and		(A, A1, A2, A3);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI31D2BWP12TLVT (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    and		(A, A1, A2, A3);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI31D4BWP12TLVT (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    and		(A, A1, A2, A3);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI32D0BWP12TLVT (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    and		(A, A1, A2, A3);
    and		(B, B1, B2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI32D1BWP12TLVT (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    and		(A, A1, A2, A3);
    and		(B, B1, B2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI32D2BWP12TLVT (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    and		(A, A1, A2, A3);
    and		(B, B1, B2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI32D4BWP12TLVT (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    and		(A, A1, A2, A3);
    and		(B, B1, B2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI32XD4BWP12TLVT (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    and		(A, A1, A2, A3);
    and		(B, B1, B2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI33D0BWP12TLVT (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    and		(A, A1, A2, A3);
    and		(B, B1, B2, B3);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI33D1BWP12TLVT (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    and		(A, A1, A2, A3);
    and		(B, B1, B2, B3);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI33D2BWP12TLVT (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    and		(A, A1, A2, A3);
    and		(B, B1, B2, B3);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI33D4BWP12TLVT (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    and		(A, A1, A2, A3);
    and		(B, B1, B2, B3);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI33XD4BWP12TLVT (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    and		(A, A1, A2, A3);
    and		(B, B1, B2, B3);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BENCD1BWP12TLVT (M0, M1, M2, X2, A, S);
    input M0, M1, M2;
    output X2, A, S;
    not          (M0N,M0);
    not          (M1N,M1);
    not          (M2N,M2);
    or           (M_temp,M0N,M1N);
    or           (M_temp1,M0,M1);
    xor          (X2N,M1,M0);
    not          (X2,X2N);
    nand         (A,M_temp1,M2N);
    nand         (S,M_temp,M2);

  specify
    (M0 => A) = (0, 0);
    (M1 => A) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b1)
    (M2 => A) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b0)
    (M2 => A) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b1)
    (M2 => A) = (0, 0);
    ifnone (M2 => A) = (0, 0);
    (M0 => S) = (0, 0);
    (M1 => S) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b0)
    (M2 => S) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b1)
    (M2 => S) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b0)
    (M2 => S) = (0, 0);
    ifnone (M2 => S) = (0, 0);
    if (M1 == 1'b1)
    (M0 => X2) = (0, 0);
    if (M1 == 1'b0)
    (M0 => X2) = (0, 0);
    ifnone (M0 => X2) = (0, 0);
    if (M0 == 1'b1)
    (M1 => X2) = (0, 0);
    if (M0 == 1'b0)
    (M1 => X2) = (0, 0);
    ifnone (M1 => X2) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BENCD2BWP12TLVT (M0, M1, M2, X2, A, S);
    input M0, M1, M2;
    output X2, A, S;
    not          (M0N,M0);
    not          (M1N,M1);
    not          (M2N,M2);
    or           (M_temp,M0N,M1N);
    or           (M_temp1,M0,M1);
    xor          (X2N,M1,M0);
    not          (X2,X2N);
    nand         (A,M_temp1,M2N);
    nand         (S,M_temp,M2);

  specify
    (M0 => A) = (0, 0);
    (M1 => A) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b1)
    (M2 => A) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b0)
    (M2 => A) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b1)
    (M2 => A) = (0, 0);
    ifnone (M2 => A) = (0, 0);
    (M0 => S) = (0, 0);
    (M1 => S) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b0)
    (M2 => S) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b1)
    (M2 => S) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b0)
    (M2 => S) = (0, 0);
    ifnone (M2 => S) = (0, 0);
    if (M1 == 1'b1)
    (M0 => X2) = (0, 0);
    if (M1 == 1'b0)
    (M0 => X2) = (0, 0);
    ifnone (M0 => X2) = (0, 0);
    if (M0 == 1'b1)
    (M1 => X2) = (0, 0);
    if (M0 == 1'b0)
    (M1 => X2) = (0, 0);
    ifnone (M1 => X2) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BENCD4BWP12TLVT (M0, M1, M2, X2, A, S);
    input M0, M1, M2;
    output X2, A, S;
    not          (M0N,M0);
    not          (M1N,M1);
    not          (M2N,M2);
    or           (M_temp,M0N,M1N);
    or           (M_temp1,M0,M1);
    xor          (X2N,M1,M0);
    not          (X2,X2N);
    nand         (A,M_temp1,M2N);
    nand         (S,M_temp,M2);

  specify
    (M0 => A) = (0, 0);
    (M1 => A) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b1)
    (M2 => A) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b0)
    (M2 => A) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b1)
    (M2 => A) = (0, 0);
    ifnone (M2 => A) = (0, 0);
    (M0 => S) = (0, 0);
    (M1 => S) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b0)
    (M2 => S) = (0, 0);
    if (M0 == 1'b0 && M1 == 1'b1)
    (M2 => S) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b0)
    (M2 => S) = (0, 0);
    ifnone (M2 => S) = (0, 0);
    if (M1 == 1'b1)
    (M0 => X2) = (0, 0);
    if (M1 == 1'b0)
    (M0 => X2) = (0, 0);
    ifnone (M0 => X2) = (0, 0);
    if (M0 == 1'b1)
    (M1 => X2) = (0, 0);
    if (M0 == 1'b0)
    (M1 => X2) = (0, 0);
    ifnone (M1 => X2) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BHDBWP12TLVT (Z);
   inout Z;
   not(weak0,weak1) (Z, Z_buf);
   not              (Z_buf, Z);

endmodule
`endcelldefine

`celldefine
module BMLD1BWP12TLVT (X2, A, S, M0, M1, PP);
   input X2, A, S, M0, M1;
   output PP;
   tsmc_mux (I0_out, S, A, M0);
   tsmc_mux (I1_out, S, A, M1);
   tsmc_mux (I2_out, I1_out, I0_out, X2);
   not (PP, I2_out);

  specify
    if (M0 == 1'b0 && M1 == 1'b1 && S == 1'b0 && X2 == 1'b0)
    (A => PP) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b1 && S == 1'b1 && X2 == 1'b1)
    (A => PP) = (0, 0);
    ifnone (A => PP) = (0, 0);
    if (A == 1'b0 && M1 == 1'b0 && S == 1'b1 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b0 && M1 == 1'b1 && S == 1'b1 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b1 && M1 == 1'b0 && S == 1'b0 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b1 && M1 == 1'b1 && S == 1'b0 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    ifnone (M0 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && S == 1'b1 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b1 && S == 1'b1 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && S == 1'b0 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b1 && S == 1'b0 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    ifnone (M1 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && M1 == 1'b0 && X2 == 1'b0)
    (S => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && M1 == 1'b1 && X2 == 1'b1)
    (S => PP) = (0, 0);
    ifnone (S => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b1 && M1 == 1'b0 && S == 1'b1)
    (X2 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && M1 == 1'b1 && S == 1'b0)
    (X2 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && M1 == 1'b1 && S == 1'b1)
    (X2 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b1 && M1 == 1'b0 && S == 1'b0)
    (X2 => PP) = (0, 0);
    ifnone (X2 => PP) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BMLD2BWP12TLVT (X2, A, S, M0, M1, PP);
   input X2, A, S, M0, M1;
   output PP;
   tsmc_mux (I0_out, S, A, M0);
   tsmc_mux (I1_out, S, A, M1);
   tsmc_mux (I2_out, I1_out, I0_out, X2);
   not (PP, I2_out);

  specify
    if (M0 == 1'b0 && M1 == 1'b1 && S == 1'b0 && X2 == 1'b0)
    (A => PP) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b1 && S == 1'b1 && X2 == 1'b1)
    (A => PP) = (0, 0);
    ifnone (A => PP) = (0, 0);
    if (A == 1'b0 && M1 == 1'b0 && S == 1'b1 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b0 && M1 == 1'b1 && S == 1'b1 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b1 && M1 == 1'b0 && S == 1'b0 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b1 && M1 == 1'b1 && S == 1'b0 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    ifnone (M0 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && S == 1'b1 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b1 && S == 1'b1 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && S == 1'b0 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b1 && S == 1'b0 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    ifnone (M1 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && M1 == 1'b0 && X2 == 1'b0)
    (S => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && M1 == 1'b1 && X2 == 1'b1)
    (S => PP) = (0, 0);
    ifnone (S => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b1 && M1 == 1'b0 && S == 1'b1)
    (X2 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && M1 == 1'b1 && S == 1'b0)
    (X2 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && M1 == 1'b1 && S == 1'b1)
    (X2 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b1 && M1 == 1'b0 && S == 1'b0)
    (X2 => PP) = (0, 0);
    ifnone (X2 => PP) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BMLD4BWP12TLVT (X2, A, S, M0, M1, PP);
   input X2, A, S, M0, M1;
   output PP;
   tsmc_mux (I0_out, S, A, M0);
   tsmc_mux (I1_out, S, A, M1);
   tsmc_mux (I2_out, I1_out, I0_out, X2);
   not (PP, I2_out);

  specify
    if (M0 == 1'b0 && M1 == 1'b1 && S == 1'b0 && X2 == 1'b0)
    (A => PP) = (0, 0);
    if (M0 == 1'b1 && M1 == 1'b1 && S == 1'b1 && X2 == 1'b1)
    (A => PP) = (0, 0);
    ifnone (A => PP) = (0, 0);
    if (A == 1'b0 && M1 == 1'b0 && S == 1'b1 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b0 && M1 == 1'b1 && S == 1'b1 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b1 && M1 == 1'b0 && S == 1'b0 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    if (A == 1'b1 && M1 == 1'b1 && S == 1'b0 && X2 == 1'b1)
    (M0 => PP) = (0, 0);
    ifnone (M0 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && S == 1'b1 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b1 && S == 1'b1 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && S == 1'b0 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b1 && S == 1'b0 && X2 == 1'b0)
    (M1 => PP) = (0, 0);
    ifnone (M1 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && M1 == 1'b0 && X2 == 1'b0)
    (S => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && M1 == 1'b1 && X2 == 1'b1)
    (S => PP) = (0, 0);
    ifnone (S => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b1 && M1 == 1'b0 && S == 1'b1)
    (X2 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b0 && M1 == 1'b1 && S == 1'b0)
    (X2 => PP) = (0, 0);
    if (A == 1'b0 && M0 == 1'b0 && M1 == 1'b1 && S == 1'b1)
    (X2 => PP) = (0, 0);
    if (A == 1'b1 && M0 == 1'b1 && M1 == 1'b0 && S == 1'b0)
    (X2 => PP) = (0, 0);
    ifnone (X2 => PP) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD0BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD12BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD16BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD1BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD20BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD24BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD2BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD3BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD4BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD6BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD8BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD0BWP12TLVT (I, OE, Z);
    input I, OE;
    output Z;
    bufif1	(Z, I, OE);
    always @(Z)
       begin
         if (!$test$plusargs("bus_conflict_off"))
            if ($countdrivers(Z) && (Z === 1'bx))
                $display("%t ++BUS CONFLICT++ : %m", $realtime);
       end

  specify
    (I => Z) = (0, 0);
    (negedge OE => (Z:I)) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD12BWP12TLVT (I, OE, Z);
    input I, OE;
    output Z;
    bufif1	(Z, I, OE);
    always @(Z)
       begin
         if (!$test$plusargs("bus_conflict_off"))
            if ($countdrivers(Z) && (Z === 1'bx))
                $display("%t ++BUS CONFLICT++ : %m", $realtime);
       end

  specify
    (I => Z) = (0, 0);
    (negedge OE => (Z:I)) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD16BWP12TLVT (I, OE, Z);
    input I, OE;
    output Z;
    bufif1	(Z, I, OE);
    always @(Z)
       begin
         if (!$test$plusargs("bus_conflict_off"))
            if ($countdrivers(Z) && (Z === 1'bx))
                $display("%t ++BUS CONFLICT++ : %m", $realtime);
       end

  specify
    (I => Z) = (0, 0);
    (negedge OE => (Z:I)) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD1BWP12TLVT (I, OE, Z);
    input I, OE;
    output Z;
    bufif1	(Z, I, OE);
    always @(Z)
       begin
         if (!$test$plusargs("bus_conflict_off"))
            if ($countdrivers(Z) && (Z === 1'bx))
                $display("%t ++BUS CONFLICT++ : %m", $realtime);
       end

  specify
    (I => Z) = (0, 0);
    (negedge OE => (Z:I)) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD20BWP12TLVT (I, OE, Z);
    input I, OE;
    output Z;
    bufif1	(Z, I, OE);
    always @(Z)
       begin
         if (!$test$plusargs("bus_conflict_off"))
            if ($countdrivers(Z) && (Z === 1'bx))
                $display("%t ++BUS CONFLICT++ : %m", $realtime);
       end

  specify
    (I => Z) = (0, 0);
    (negedge OE => (Z:I)) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD24BWP12TLVT (I, OE, Z);
    input I, OE;
    output Z;
    bufif1	(Z, I, OE);
    always @(Z)
       begin
         if (!$test$plusargs("bus_conflict_off"))
            if ($countdrivers(Z) && (Z === 1'bx))
                $display("%t ++BUS CONFLICT++ : %m", $realtime);
       end

  specify
    (I => Z) = (0, 0);
    (negedge OE => (Z:I)) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD2BWP12TLVT (I, OE, Z);
    input I, OE;
    output Z;
    bufif1	(Z, I, OE);
    always @(Z)
       begin
         if (!$test$plusargs("bus_conflict_off"))
            if ($countdrivers(Z) && (Z === 1'bx))
                $display("%t ++BUS CONFLICT++ : %m", $realtime);
       end

  specify
    (I => Z) = (0, 0);
    (negedge OE => (Z:I)) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD3BWP12TLVT (I, OE, Z);
    input I, OE;
    output Z;
    bufif1	(Z, I, OE);
    always @(Z)
       begin
         if (!$test$plusargs("bus_conflict_off"))
            if ($countdrivers(Z) && (Z === 1'bx))
                $display("%t ++BUS CONFLICT++ : %m", $realtime);
       end

  specify
    (I => Z) = (0, 0);
    (negedge OE => (Z:I)) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD4BWP12TLVT (I, OE, Z);
    input I, OE;
    output Z;
    bufif1	(Z, I, OE);
    always @(Z)
       begin
         if (!$test$plusargs("bus_conflict_off"))
            if ($countdrivers(Z) && (Z === 1'bx))
                $display("%t ++BUS CONFLICT++ : %m", $realtime);
       end

  specify
    (I => Z) = (0, 0);
    (negedge OE => (Z:I)) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD6BWP12TLVT (I, OE, Z);
    input I, OE;
    output Z;
    bufif1	(Z, I, OE);
    always @(Z)
       begin
         if (!$test$plusargs("bus_conflict_off"))
            if ($countdrivers(Z) && (Z === 1'bx))
                $display("%t ++BUS CONFLICT++ : %m", $realtime);
       end

  specify
    (I => Z) = (0, 0);
    (negedge OE => (Z:I)) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD8BWP12TLVT (I, OE, Z);
    input I, OE;
    output Z;
    bufif1	(Z, I, OE);
    always @(Z)
       begin
         if (!$test$plusargs("bus_conflict_off"))
            if ($countdrivers(Z) && (Z === 1'bx))
                $display("%t ++BUS CONFLICT++ : %m", $realtime);
       end

  specify
    (I => Z) = (0, 0);
    (negedge OE => (Z:I)) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKAN2D0BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKAN2D1BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKAN2D2BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKAN2D4BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKAN2D8BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD0BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD12BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD16BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD1BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD20BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD24BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD2BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD3BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD4BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD6BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD8BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKLHQD12BWP12TLVT ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    // Dummy Buffer
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, CPN_d, E_d ;
    buf ( _TE, TE_d );
    buf ( _CPN, CPN_d );
    buf ( _E, E_d );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `else 	// Reserve for non NTC.
    buf ( _TE, TE );
    buf ( _CPN, CPN );
    buf ( _E, E );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CPN => Q) = (0, 0);
    $width (posedge CPN, 0, 0, notifier);
    $width (negedge CPN, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD16BWP12TLVT ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    // Dummy Buffer
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, CPN_d, E_d ;
    buf ( _TE, TE_d );
    buf ( _CPN, CPN_d );
    buf ( _E, E_d );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `else 	// Reserve for non NTC.
    buf ( _TE, TE );
    buf ( _CPN, CPN );
    buf ( _E, E );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CPN => Q) = (0, 0);
    $width (posedge CPN, 0, 0, notifier);
    $width (negedge CPN, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD1BWP12TLVT ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    // Dummy Buffer
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, CPN_d, E_d ;
    buf ( _TE, TE_d );
    buf ( _CPN, CPN_d );
    buf ( _E, E_d );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `else 	// Reserve for non NTC.
    buf ( _TE, TE );
    buf ( _CPN, CPN );
    buf ( _E, E );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CPN => Q) = (0, 0);
    $width (posedge CPN, 0, 0, notifier);
    $width (negedge CPN, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD20BWP12TLVT ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    // Dummy Buffer
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, CPN_d, E_d ;
    buf ( _TE, TE_d );
    buf ( _CPN, CPN_d );
    buf ( _E, E_d );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `else 	// Reserve for non NTC.
    buf ( _TE, TE );
    buf ( _CPN, CPN );
    buf ( _E, E );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CPN => Q) = (0, 0);
    $width (posedge CPN, 0, 0, notifier);
    $width (negedge CPN, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD24BWP12TLVT ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    // Dummy Buffer
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, CPN_d, E_d ;
    buf ( _TE, TE_d );
    buf ( _CPN, CPN_d );
    buf ( _E, E_d );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `else 	// Reserve for non NTC.
    buf ( _TE, TE );
    buf ( _CPN, CPN );
    buf ( _E, E );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CPN => Q) = (0, 0);
    $width (posedge CPN, 0, 0, notifier);
    $width (negedge CPN, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD2BWP12TLVT ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    // Dummy Buffer
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, CPN_d, E_d ;
    buf ( _TE, TE_d );
    buf ( _CPN, CPN_d );
    buf ( _E, E_d );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `else 	// Reserve for non NTC.
    buf ( _TE, TE );
    buf ( _CPN, CPN );
    buf ( _E, E );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CPN => Q) = (0, 0);
    $width (posedge CPN, 0, 0, notifier);
    $width (negedge CPN, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD3BWP12TLVT ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    // Dummy Buffer
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, CPN_d, E_d ;
    buf ( _TE, TE_d );
    buf ( _CPN, CPN_d );
    buf ( _E, E_d );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `else 	// Reserve for non NTC.
    buf ( _TE, TE );
    buf ( _CPN, CPN );
    buf ( _E, E );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CPN => Q) = (0, 0);
    $width (posedge CPN, 0, 0, notifier);
    $width (negedge CPN, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD4BWP12TLVT ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    // Dummy Buffer
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, CPN_d, E_d ;
    buf ( _TE, TE_d );
    buf ( _CPN, CPN_d );
    buf ( _E, E_d );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `else 	// Reserve for non NTC.
    buf ( _TE, TE );
    buf ( _CPN, CPN );
    buf ( _E, E );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CPN => Q) = (0, 0);
    $width (posedge CPN, 0, 0, notifier);
    $width (negedge CPN, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD6BWP12TLVT ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    // Dummy Buffer
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, CPN_d, E_d ;
    buf ( _TE, TE_d );
    buf ( _CPN, CPN_d );
    buf ( _E, E_d );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `else 	// Reserve for non NTC.
    buf ( _TE, TE );
    buf ( _CPN, CPN );
    buf ( _E, E );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CPN => Q) = (0, 0);
    $width (posedge CPN, 0, 0, notifier);
    $width (negedge CPN, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD8BWP12TLVT ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    // Dummy Buffer
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, CPN_d, E_d ;
    buf ( _TE, TE_d );
    buf ( _CPN, CPN_d );
    buf ( _E, E_d );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `else 	// Reserve for non NTC.
    buf ( _TE, TE );
    buf ( _CPN, CPN );
    buf ( _E, E );
    or ( _G001, _E, _TE );
    tsmc_dla ( _enl, _G001, _CPN, 1'b1, 1'b1, notifier );
    not ( _enlb, _enl );
    or ( Q, _enlb, _CPN );
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CPN => Q) = (0, 0);
    $width (posedge CPN, 0, 0, notifier);
    $width (negedge CPN, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (negedge CPN &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD12BWP12TLVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, E_d, CP_d ;
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E_d, TE_d);
    not		(CPB, CP_d);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP_d);
  `else 	// Reserve for non NTC.
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E, TE);
    not		(CPB, CP);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CP => Q) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD16BWP12TLVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, E_d, CP_d ;
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E_d, TE_d);
    not		(CPB, CP_d);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP_d);
  `else 	// Reserve for non NTC.
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E, TE);
    not		(CPB, CP);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CP => Q) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD1BWP12TLVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, E_d, CP_d ;
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E_d, TE_d);
    not		(CPB, CP_d);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP_d);
  `else 	// Reserve for non NTC.
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E, TE);
    not		(CPB, CP);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CP => Q) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD20BWP12TLVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, E_d, CP_d ;
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E_d, TE_d);
    not		(CPB, CP_d);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP_d);
  `else 	// Reserve for non NTC.
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E, TE);
    not		(CPB, CP);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CP => Q) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD24BWP12TLVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, E_d, CP_d ;
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E_d, TE_d);
    not		(CPB, CP_d);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP_d);
  `else 	// Reserve for non NTC.
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E, TE);
    not		(CPB, CP);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CP => Q) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD2BWP12TLVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, E_d, CP_d ;
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E_d, TE_d);
    not		(CPB, CP_d);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP_d);
  `else 	// Reserve for non NTC.
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E, TE);
    not		(CPB, CP);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CP => Q) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD3BWP12TLVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, E_d, CP_d ;
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E_d, TE_d);
    not		(CPB, CP_d);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP_d);
  `else 	// Reserve for non NTC.
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E, TE);
    not		(CPB, CP);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CP => Q) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD4BWP12TLVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, E_d, CP_d ;
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E_d, TE_d);
    not		(CPB, CP_d);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP_d);
  `else 	// Reserve for non NTC.
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E, TE);
    not		(CPB, CP);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CP => Q) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD6BWP12TLVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, E_d, CP_d ;
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E_d, TE_d);
    not		(CPB, CP_d);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP_d);
  `else 	// Reserve for non NTC.
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E, TE);
    not		(CPB, CP);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CP => Q) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD8BWP12TLVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire TE_d, E_d, CP_d ;
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E_d, TE_d);
    not		(CPB, CP_d);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP_d);
  `else 	// Reserve for non NTC.
    pullup	(CDN);
    pullup	(SDN);
    or		(D_i, E, TE);
    not		(CPB, CP);
    tsmc_dla 	(Q_buf, D_i, CPB, CDN, SDN, notifier);
    and         (Q, Q_buf, CP);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (TE_int_not, TE_d);
  `else
    not  (E_int_not, E);
    not  (TE_int_not, TE);
  `endif
    buf  (E_check, TE_int_not);
  buf  (TE_check, E_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CP => Q) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, posedge TE, 0, 0, notifier);
    $setuphold (posedge CP &&& TE_DEFCHK, negedge TE, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKMUX2D0BWP12TLVT (I0, I1, S, Z);
   input I0, I1, S;
   output Z;
   tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    ifnone (I0 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    ifnone (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
    ifnone (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKMUX2D1BWP12TLVT (I0, I1, S, Z);
   input I0, I1, S;
   output Z;
   tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    ifnone (I0 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    ifnone (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
    ifnone (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKMUX2D2BWP12TLVT (I0, I1, S, Z);
   input I0, I1, S;
   output Z;
   tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    ifnone (I0 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    ifnone (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
    ifnone (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKMUX2D4BWP12TLVT (I0, I1, S, Z);
   input I0, I1, S;
   output Z;
   tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    ifnone (I0 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    ifnone (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
    ifnone (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND0BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND12BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND16BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND1BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND20BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND24BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2D0BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nand		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2D1BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nand		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2D2BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nand		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2D3BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nand		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2D4BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nand		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2D8BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nand		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND3BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND4BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND6BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND8BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKXOR2D0BWP12TLVT (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
  xor		(Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    ifnone (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
    ifnone (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKXOR2D1BWP12TLVT (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
  xor		(Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    ifnone (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
    ifnone (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKXOR2D2BWP12TLVT (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
  xor		(Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    ifnone (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
    ifnone (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKXOR2D4BWP12TLVT (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
  xor		(Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    ifnone (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
    ifnone (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CMPE42D1BWP12TLVT (A, B, C, D, CIX, S, COX, CO);
input A, B, C, D, CIX;
output S, COX, CO;
  xor  (temp1, A, B);
  xor  (IS, temp1, C);
  and  (temp2, A, B);
  and  (temp3, A, C);
  and  (temp5, B, C);
  or   (COX, temp2, temp3, temp5);
  xor  (temp6, IS, D);
  xor  (S, temp6, CIX);
  and  (temp7, IS, D);
  and  (temp8, IS, CIX);
  and  (temp9, D, CIX);
  or   (CO, temp7, temp8, temp9);

  specify
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (A => CO) = (0, 0);
    ifnone (A => CO) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (B => CO) = (0, 0);
    ifnone (B => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (C => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (C => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (C => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (C => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (C => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (C => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (C => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (C => CO) = (0, 0);
    ifnone (C => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b1)
    (CIX => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0)
    (CIX => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0)
    (CIX => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b1)
    (CIX => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0)
    (CIX => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1)
    (CIX => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1)
    (CIX => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0)
    (CIX => CO) = (0, 0);
    ifnone (CIX => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && CIX == 1'b1)
    (D => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && CIX == 1'b0)
    (D => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && CIX == 1'b0)
    (D => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && CIX == 1'b1)
    (D => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && CIX == 1'b0)
    (D => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && CIX == 1'b1)
    (D => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && CIX == 1'b1)
    (D => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && CIX == 1'b0)
    (D => CO) = (0, 0);
    ifnone (D => CO) = (0, 0);
    if (B == 1'b0 && C == 1'b1)
    (A => COX) = (0, 0);
    if (B == 1'b1 && C == 1'b0)
    (A => COX) = (0, 0);
    ifnone (A => COX) = (0, 0);
    if (A == 1'b0 && C == 1'b1)
    (B => COX) = (0, 0);
    if (A == 1'b1 && C == 1'b0)
    (B => COX) = (0, 0);
    ifnone (B => COX) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (C => COX) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (C => COX) = (0, 0);
    ifnone (C => COX) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (C => S) = (0, 0);
    ifnone (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0)
    (CIX => S) = (0, 0);
    ifnone (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && CIX == 1'b0)
    (D => S) = (0, 0);
    ifnone (D => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CMPE42D2BWP12TLVT (A, B, C, D, CIX, S, COX, CO);
input A, B, C, D, CIX;
output S, COX, CO;
  xor  (temp1, A, B);
  xor  (IS, temp1, C);
  and  (temp2, A, B);
  and  (temp3, A, C);
  and  (temp5, B, C);
  or   (COX, temp2, temp3, temp5);
  xor  (temp6, IS, D);
  xor  (S, temp6, CIX);
  and  (temp7, IS, D);
  and  (temp8, IS, CIX);
  and  (temp9, D, CIX);
  or   (CO, temp7, temp8, temp9);

  specify
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (A => CO) = (0, 0);
    ifnone (A => CO) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (B => CO) = (0, 0);
    ifnone (B => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (C => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (C => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (C => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (C => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (C => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (C => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (C => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (C => CO) = (0, 0);
    ifnone (C => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b1)
    (CIX => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0)
    (CIX => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0)
    (CIX => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b1)
    (CIX => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0)
    (CIX => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1)
    (CIX => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1)
    (CIX => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0)
    (CIX => CO) = (0, 0);
    ifnone (CIX => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && CIX == 1'b1)
    (D => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && CIX == 1'b0)
    (D => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && CIX == 1'b0)
    (D => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && CIX == 1'b1)
    (D => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && CIX == 1'b0)
    (D => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && CIX == 1'b1)
    (D => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && CIX == 1'b1)
    (D => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && CIX == 1'b0)
    (D => CO) = (0, 0);
    ifnone (D => CO) = (0, 0);
    if (B == 1'b0 && C == 1'b1)
    (A => COX) = (0, 0);
    if (B == 1'b1 && C == 1'b0)
    (A => COX) = (0, 0);
    ifnone (A => COX) = (0, 0);
    if (A == 1'b0 && C == 1'b1)
    (B => COX) = (0, 0);
    if (A == 1'b1 && C == 1'b0)
    (B => COX) = (0, 0);
    ifnone (B => COX) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (C => COX) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (C => COX) = (0, 0);
    ifnone (C => COX) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b0 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIX == 1'b1 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b0 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIX == 1'b1 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b0 && D == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIX == 1'b1 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b0 && D == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIX == 1'b1 && D == 1'b0)
    (C => S) = (0, 0);
    ifnone (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && D == 1'b0)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && D == 1'b1)
    (CIX => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && D == 1'b0)
    (CIX => S) = (0, 0);
    ifnone (CIX => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b0 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && C == 1'b1 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b0 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && C == 1'b1 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b0 && CIX == 1'b0)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && C == 1'b1 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b0 && CIX == 1'b1)
    (D => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && C == 1'b1 && CIX == 1'b0)
    (D => S) = (0, 0);
    ifnone (D => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DCAP16BWP12TLVT;
    // No function
endmodule
`endcelldefine

`celldefine
module DCAP32BWP12TLVT;
    // No function
endmodule
`endcelldefine

`celldefine
module DCAP4BWP12TLVT;
    // No function
endmodule
`endcelldefine

`celldefine
module DCAP64BWP12TLVT;
    // No function
endmodule
`endcelldefine

`celldefine
module DCAP8BWP12TLVT;
    // No function
endmodule
`endcelldefine

`celldefine
module DCAPBWP12TLVT;
    // No function
endmodule
`endcelldefine

`celldefine
module DEL005BWP12TLVT (I, Z);
    input I;
    output Z;
    buf         (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL015BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL01BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL02BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL0BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL1BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL2BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL3BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL4BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DFCND1BWP12TLVT (D, CP, CDN, Q, QN);
    input D, CP, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire D_d, CP_d ;
    pullup	 (SDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    pullup	 (SDN);
    tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (CP_check, CDN_i);
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCND2BWP12TLVT (D, CP, CDN, Q, QN);
    input D, CP, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire D_d, CP_d ;
    pullup	 (SDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    pullup	 (SDN);
    tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (CP_check, CDN_i);
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCND4BWP12TLVT (D, CP, CDN, Q, QN);
    input D, CP, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire D_d, CP_d ;
    pullup	 (SDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    pullup	 (SDN);
    tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (CP_check, CDN_i);
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCNQD1BWP12TLVT (D, CP, CDN, Q);
    input D, CP, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire D_d, CP_d ;
    pullup   (SDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    pullup   (SDN);
    tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (CP_check, CDN_i);
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCNQD2BWP12TLVT (D, CP, CDN, Q);
    input D, CP, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire D_d, CP_d ;
    pullup   (SDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    pullup   (SDN);
    tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (CP_check, CDN_i);
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCNQD4BWP12TLVT (D, CP, CDN, Q);
    input D, CP, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire D_d, CP_d ;
    pullup   (SDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    pullup   (SDN);
    tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (CP_check, CDN_i);
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCSND1BWP12TLVT (D, CP, CDN, SDN, Q, QN);
    input D, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire D_d, CP_d ;
    tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (CP_check, CDN_i, SDN_i);
  and  (D_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCSND2BWP12TLVT (D, CP, CDN, SDN, Q, QN);
    input D, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire D_d, CP_d ;
    tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (CP_check, CDN_i, SDN_i);
  and  (D_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCSND4BWP12TLVT (D, CP, CDN, SDN, Q, QN);
    input D, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire D_d, CP_d ;
    tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (CP_check, CDN_i, SDN_i);
  and  (D_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCSNQD1BWP12TLVT (D, CP, CDN, SDN, Q);
    input D, CP, CDN, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire D_d, CP_d ;
    tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (CP_check, CDN_i, SDN_i);
  and  (D_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCSNQD2BWP12TLVT (D, CP, CDN, SDN, Q);
    input D, CP, CDN, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire D_d, CP_d ;
    tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (CP_check, CDN_i, SDN_i);
  and  (D_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCSNQD4BWP12TLVT (D, CP, CDN, SDN, Q);
    input D, CP, CDN, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire D_d, CP_d ;
    tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (CP_check, CDN_i, SDN_i);
  and  (D_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFD1BWP12TLVT (D, CP, Q, QN);
    input D, CP;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CP_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not	     (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not	     (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  pullup  (CP_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFD2BWP12TLVT (D, CP, Q, QN);
    input D, CP;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CP_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not	     (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not	     (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  pullup  (CP_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFD4BWP12TLVT (D, CP, Q, QN);
    input D, CP;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CP_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not	     (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not	     (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  pullup  (CP_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCND1BWP12TLVT (D, CP, CN, Q, QN);
    input D, CP, CN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CP_d, CN_d ;
    pullup   (CDN);
    pullup   (SDN);
    and      (D_i, CN_d, D_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    and      (D_i, CN, D);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (D_check, CN_d);
  `else
    buf  (D_check, CN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && D)))) = (0, 0);
    (posedge CP => (QN-:((CN && D)))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCND2BWP12TLVT (D, CP, CN, Q, QN);
    input D, CP, CN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CP_d, CN_d ;
    pullup   (CDN);
    pullup   (SDN);
    and      (D_i, CN_d, D_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    and      (D_i, CN, D);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (D_check, CN_d);
  `else
    buf  (D_check, CN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && D)))) = (0, 0);
    (posedge CP => (QN-:((CN && D)))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCND4BWP12TLVT (D, CP, CN, Q, QN);
    input D, CP, CN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CP_d, CN_d ;
    pullup   (CDN);
    pullup   (SDN);
    and      (D_i, CN_d, D_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    and      (D_i, CN, D);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (D_check, CN_d);
  `else
    buf  (D_check, CN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && D)))) = (0, 0);
    (posedge CP => (QN-:((CN && D)))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCNQD1BWP12TLVT (D, CP, CN, Q);
    input D, CP, CN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CP_d, CN_d ;
    pullup   (CDN); 
    pullup   (SDN);     
    and      (D_i, CN_d, D_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
  `else 	// Reserve for non NTC.
    pullup   (CDN); 
    pullup   (SDN);     
    and      (D_i, CN, D);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (D_check, CN_d);
  `else
    buf  (D_check, CN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && D)))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCNQD2BWP12TLVT (D, CP, CN, Q);
    input D, CP, CN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CP_d, CN_d ;
    pullup   (CDN); 
    pullup   (SDN);     
    and      (D_i, CN_d, D_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
  `else 	// Reserve for non NTC.
    pullup   (CDN); 
    pullup   (SDN);     
    and      (D_i, CN, D);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (D_check, CN_d);
  `else
    buf  (D_check, CN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && D)))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCNQD4BWP12TLVT (D, CP, CN, Q);
    input D, CP, CN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CP_d, CN_d ;
    pullup   (CDN); 
    pullup   (SDN);     
    and      (D_i, CN_d, D_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
  `else 	// Reserve for non NTC.
    pullup   (CDN); 
    pullup   (SDN);     
    and      (D_i, CN, D);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (D_check, CN_d);
  `else
    buf  (D_check, CN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && D)))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCSND1BWP12TLVT (D, CP, CN, SN, Q, QN);
    input D, CP, CN, SN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CP_d, CN_d, SN_d ;
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN_d);
    or       (DS, S, D_d);   
    and      (D_i, CN_d, DS);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN);
    or       (DS, S, D);   
    and      (D_i, CN, DS);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (SN_check, CN_d);
    and  (D_check, SN_d, CN_d);
  `else
    buf  (SN_check, CN);
    and  (D_check, SN, CN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && D) || (CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((CN && D) || (CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCSND2BWP12TLVT (D, CP, CN, SN, Q, QN);
    input D, CP, CN, SN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CP_d, CN_d, SN_d ;
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN_d);
    or       (DS, S, D_d);   
    and      (D_i, CN_d, DS);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN);
    or       (DS, S, D);   
    and      (D_i, CN, DS);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (SN_check, CN_d);
    and  (D_check, SN_d, CN_d);
  `else
    buf  (SN_check, CN);
    and  (D_check, SN, CN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && D) || (CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((CN && D) || (CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCSND4BWP12TLVT (D, CP, CN, SN, Q, QN);
    input D, CP, CN, SN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CP_d, CN_d, SN_d ;
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN_d);
    or       (DS, S, D_d);   
    and      (D_i, CN_d, DS);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN);
    or       (DS, S, D);   
    and      (D_i, CN, DS);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (SN_check, CN_d);
    and  (D_check, SN_d, CN_d);
  `else
    buf  (SN_check, CN);
    and  (D_check, SN, CN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && D) || (CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((CN && D) || (CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKSND1BWP12TLVT (D, CP, SN, Q, QN);
    input D, CP, SN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CP_d, SN_d ;
    pullup   (CDN);
    pullup   (SDN);
    not      (S, SN_d);
    or       (D_i, S, D_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    not      (S, SN);
    or       (D_i, S, D);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (D_check, SN_d);
  `else
    buf  (D_check, SN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((D) || (!(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((D) || (!(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKSND2BWP12TLVT (D, CP, SN, Q, QN);
    input D, CP, SN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CP_d, SN_d ;
    pullup   (CDN);
    pullup   (SDN);
    not      (S, SN_d);
    or       (D_i, S, D_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    not      (S, SN);
    or       (D_i, S, D);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (D_check, SN_d);
  `else
    buf  (D_check, SN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((D) || (!(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((D) || (!(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKSND4BWP12TLVT (D, CP, SN, Q, QN);
    input D, CP, SN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CP_d, SN_d ;
    pullup   (CDN);
    pullup   (SDN);
    not      (S, SN_d);
    or       (D_i, S, D_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    not      (S, SN);
    or       (D_i, S, D);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    buf  (D_check, SN_d);
  `else
    buf  (D_check, SN);
  `endif
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((D) || (!(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((D) || (!(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNCND1BWP12TLVT (D, CPN, CDN, Q, QN);
    input D, CPN, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, CPN_d ;
    pullup	(SDN);
    not		(CP, CPN_d);
    tsmc_dff	(Q_buf, D_d, CP, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup	(SDN);
    not		(CP, CPN);
    tsmc_dff	(Q_buf, D, CP, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (CPN_check, CDN_i);
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:D)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge CDN, negedge CPN, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge CDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNCND2BWP12TLVT (D, CPN, CDN, Q, QN);
    input D, CPN, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, CPN_d ;
    pullup	(SDN);
    not		(CP, CPN_d);
    tsmc_dff	(Q_buf, D_d, CP, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup	(SDN);
    not		(CP, CPN);
    tsmc_dff	(Q_buf, D, CP, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (CPN_check, CDN_i);
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:D)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge CDN, negedge CPN, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge CDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNCND4BWP12TLVT (D, CPN, CDN, Q, QN);
    input D, CPN, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, CPN_d ;
    pullup	(SDN);
    not		(CP, CPN_d);
    tsmc_dff	(Q_buf, D_d, CP, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup	(SDN);
    not		(CP, CPN);
    tsmc_dff	(Q_buf, D, CP, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (CPN_check, CDN_i);
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:D)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge CDN, negedge CPN, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge CDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNCSND1BWP12TLVT (D, CPN, CDN, SDN, Q, QN);
    input D, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf          (CDN_i, CDN_d);
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
      buf          (SDN_i, SDN);
    `endif
    wire D_d, CPN_d ;
    not		 (CP, CPN_d);
    tsmc_dff	 (Q_buf, D_d, CP, CDN_i, SDN_i, notifier);
    buf          (Q, Q_buf);
    not          (QN_buf, Q_buf);
    and          (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    buf          (SDN_i, SDN);
    not		 (CP, CPN);
    tsmc_dff	 (Q_buf, D, CP, CDN_i, SDN_i, notifier);
    buf          (Q, Q_buf);
    not          (QN_buf, Q_buf);
    and          (QN, QN_buf, SDN_i);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (CPN_check, CDN_i, SDN_i);
  and  (D_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:D)) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge CDN, negedge CPN, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, negedge CPN, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge CDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNCSND2BWP12TLVT (D, CPN, CDN, SDN, Q, QN);
    input D, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf          (CDN_i, CDN_d);
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
      buf          (SDN_i, SDN);
    `endif
    wire D_d, CPN_d ;
    not		 (CP, CPN_d);
    tsmc_dff	 (Q_buf, D_d, CP, CDN_i, SDN_i, notifier);
    buf          (Q, Q_buf);
    not          (QN_buf, Q_buf);
    and          (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    buf          (SDN_i, SDN);
    not		 (CP, CPN);
    tsmc_dff	 (Q_buf, D, CP, CDN_i, SDN_i, notifier);
    buf          (Q, Q_buf);
    not          (QN_buf, Q_buf);
    and          (QN, QN_buf, SDN_i);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (CPN_check, CDN_i, SDN_i);
  and  (D_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:D)) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge CDN, negedge CPN, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, negedge CPN, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge CDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNCSND4BWP12TLVT (D, CPN, CDN, SDN, Q, QN);
    input D, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf          (CDN_i, CDN_d);
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
      buf          (SDN_i, SDN);
    `endif
    wire D_d, CPN_d ;
    not		 (CP, CPN_d);
    tsmc_dff	 (Q_buf, D_d, CP, CDN_i, SDN_i, notifier);
    buf          (Q, Q_buf);
    not          (QN_buf, Q_buf);
    and          (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    buf          (SDN_i, SDN);
    not		 (CP, CPN);
    tsmc_dff	 (Q_buf, D, CP, CDN_i, SDN_i, notifier);
    buf          (Q, Q_buf);
    not          (QN_buf, Q_buf);
    and          (QN, QN_buf, SDN_i);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (CPN_check, CDN_i, SDN_i);
  and  (D_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:D)) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge CDN, negedge CPN, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, negedge CPN, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge CDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFND1BWP12TLVT (D, CPN, Q, QN);
    input D, CPN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CPN_d ;
    pullup	(CDN);
    pullup      (SDN);
    not		(CP, CPN_d);
    tsmc_dff	(Q_buf, D_d, CP, CDN, SDN, notifier);
    buf         (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup	(CDN);
    pullup      (SDN);
    not		(CP, CPN);
    tsmc_dff	(Q_buf, D, CP, CDN, SDN, notifier);
    buf         (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  pullup  (CPN_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:D)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFND2BWP12TLVT (D, CPN, Q, QN);
    input D, CPN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CPN_d ;
    pullup	(CDN);
    pullup      (SDN);
    not		(CP, CPN_d);
    tsmc_dff	(Q_buf, D_d, CP, CDN, SDN, notifier);
    buf         (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup	(CDN);
    pullup      (SDN);
    not		(CP, CPN);
    tsmc_dff	(Q_buf, D, CP, CDN, SDN, notifier);
    buf         (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  pullup  (CPN_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:D)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFND4BWP12TLVT (D, CPN, Q, QN);
    input D, CPN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CPN_d ;
    pullup	(CDN);
    pullup      (SDN);
    not		(CP, CPN_d);
    tsmc_dff	(Q_buf, D_d, CP, CDN, SDN, notifier);
    buf         (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup	(CDN);
    pullup      (SDN);
    not		(CP, CPN);
    tsmc_dff	(Q_buf, D, CP, CDN, SDN, notifier);
    buf         (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  pullup  (CPN_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:D)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNSND1BWP12TLVT (D, CPN, SDN, Q, QN);
    input D, CPN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, CPN_d ;
    pullup	(CDN);
    not		(CP, CPN_d);
    tsmc_dff	(Q_buf, D_d, CP, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup	(CDN);
    not		(CP, CPN);
    tsmc_dff	(Q_buf, D, CP, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (CPN_check, SDN_i);
  buf  (D_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:D)) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge SDN, negedge CPN, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge SDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNSND2BWP12TLVT (D, CPN, SDN, Q, QN);
    input D, CPN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, CPN_d ;
    pullup	(CDN);
    not		(CP, CPN_d);
    tsmc_dff	(Q_buf, D_d, CP, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup	(CDN);
    not		(CP, CPN);
    tsmc_dff	(Q_buf, D, CP, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (CPN_check, SDN_i);
  buf  (D_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:D)) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge SDN, negedge CPN, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge SDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNSND4BWP12TLVT (D, CPN, SDN, Q, QN);
    input D, CPN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, CPN_d ;
    pullup	(CDN);
    not		(CP, CPN_d);
    tsmc_dff	(Q_buf, D_d, CP, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup	(CDN);
    not		(CP, CPN);
    tsmc_dff	(Q_buf, D, CP, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (CPN_check, SDN_i);
  buf  (D_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:D)) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge SDN, negedge CPN, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge SDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFQD1BWP12TLVT (D, CP, Q);
    input D, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CP_d ;
    pullup	 (CDN);
    pullup	 (SDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup	 (CDN);
    pullup	 (SDN);
    tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  pullup  (CP_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFQD2BWP12TLVT (D, CP, Q);
    input D, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CP_d ;
    pullup	 (CDN);
    pullup	 (SDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup	 (CDN);
    pullup	 (SDN);
    tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  pullup  (CP_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFQD4BWP12TLVT (D, CP, Q);
    input D, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CP_d ;
    pullup	 (CDN);
    pullup	 (SDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup	 (CDN);
    pullup	 (SDN);
    tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  pullup  (CP_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFSND1BWP12TLVT (D, CP, SDN, Q, QN);
    input D, CP, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (SDN_i, SDN);
    `endif
    wire D_d, CP_d ;
    pullup   (CDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (SDN_i, SDN);
    pullup   (CDN);
    tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (CP_check, SDN_i);
  buf  (D_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFSND2BWP12TLVT (D, CP, SDN, Q, QN);
    input D, CP, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (SDN_i, SDN);
    `endif
    wire D_d, CP_d ;
    pullup   (CDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (SDN_i, SDN);
    pullup   (CDN);
    tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (CP_check, SDN_i);
  buf  (D_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFSND4BWP12TLVT (D, CP, SDN, Q, QN);
    input D, CP, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (SDN_i, SDN);
    `endif
    wire D_d, CP_d ;
    pullup   (CDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (SDN_i, SDN);
    pullup   (CDN);
    tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (CP_check, SDN_i);
  buf  (D_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFSNQD1BWP12TLVT (D, CP, SDN, Q);
    input D, CP, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (SDN_i, SDN);
    `endif
    wire D_d, CP_d ;
    pullup   (CDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (SDN_i, SDN);
    pullup   (CDN);
    tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (CP_check, SDN_i);
  buf  (D_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFSNQD2BWP12TLVT (D, CP, SDN, Q);
    input D, CP, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (SDN_i, SDN);
    `endif
    wire D_d, CP_d ;
    pullup   (CDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (SDN_i, SDN);
    pullup   (CDN);
    tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (CP_check, SDN_i);
  buf  (D_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFSNQD4BWP12TLVT (D, CP, SDN, Q);
    input D, CP, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (SDN_i, SDN);
    `endif
    wire D_d, CP_d ;
    pullup   (CDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (SDN_i, SDN);
    pullup   (CDN);
    tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (CP_check, SDN_i);
  buf  (D_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFXD1BWP12TLVT (DA, DB, SA, CP, Q, QN);
    input DA, DB, SA, CP;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire DA_d, DB_d, SA_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB_d, DA_d, SA_d);
    tsmc_dff     (Q_buf, D, CP_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB, DA, SA);
    tsmc_dff     (Q_buf, D, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    buf  (DA_check, SA_d);
  `else
    not  (SA_int_not, SA);
    buf  (DA_check, SA);
  `endif
  buf  (DB_check, SA_int_not);
  pullup  (CP_check);
  pullup  (SA_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    (posedge CP => (QN-:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier,,, CP_d, SA_d);
  `else
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFXD2BWP12TLVT (DA, DB, SA, CP, Q, QN);
    input DA, DB, SA, CP;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire DA_d, DB_d, SA_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB_d, DA_d, SA_d);
    tsmc_dff     (Q_buf, D, CP_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB, DA, SA);
    tsmc_dff     (Q_buf, D, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    buf  (DA_check, SA_d);
  `else
    not  (SA_int_not, SA);
    buf  (DA_check, SA);
  `endif
  buf  (DB_check, SA_int_not);
  pullup  (CP_check);
  pullup  (SA_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    (posedge CP => (QN-:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier,,, CP_d, SA_d);
  `else
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFXD4BWP12TLVT (DA, DB, SA, CP, Q, QN);
    input DA, DB, SA, CP;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire DA_d, DB_d, SA_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB_d, DA_d, SA_d);
    tsmc_dff     (Q_buf, D, CP_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB, DA, SA);
    tsmc_dff     (Q_buf, D, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    buf  (DA_check, SA_d);
  `else
    not  (SA_int_not, SA);
    buf  (DA_check, SA);
  `endif
  buf  (DB_check, SA_int_not);
  pullup  (CP_check);
  pullup  (SA_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    (posedge CP => (QN-:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier,,, CP_d, SA_d);
  `else
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFXQD1BWP12TLVT (DA, DB, SA, CP, Q);
    input DA, DB, SA, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire DA_d, DB_d, SA_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB_d, DA_d, SA_d);
    tsmc_dff     (Q_buf, D, CP_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB, DA, SA);
    tsmc_dff     (Q_buf, D, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    buf  (DA_check, SA_d);
  `else
    not  (SA_int_not, SA);
    buf  (DA_check, SA);
  `endif
  buf  (DB_check, SA_int_not);
  pullup  (CP_check);
  pullup  (SA_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier,,, CP_d, SA_d);
  `else
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFXQD2BWP12TLVT (DA, DB, SA, CP, Q);
    input DA, DB, SA, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire DA_d, DB_d, SA_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB_d, DA_d, SA_d);
    tsmc_dff     (Q_buf, D, CP_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB, DA, SA);
    tsmc_dff     (Q_buf, D, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    buf  (DA_check, SA_d);
  `else
    not  (SA_int_not, SA);
    buf  (DA_check, SA);
  `endif
  buf  (DB_check, SA_int_not);
  pullup  (CP_check);
  pullup  (SA_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier,,, CP_d, SA_d);
  `else
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFXQD4BWP12TLVT (DA, DB, SA, CP, Q);
    input DA, DB, SA, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire DA_d, DB_d, SA_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB_d, DA_d, SA_d);
    tsmc_dff     (Q_buf, D, CP_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB, DA, SA);
    tsmc_dff     (Q_buf, D, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    buf  (DA_check, SA_d);
  `else
    not  (SA_int_not, SA);
    buf  (DA_check, SA);
  `endif
  buf  (DB_check, SA_int_not);
  pullup  (CP_check);
  pullup  (SA_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier,,, CP_d, SA_d);
  `else
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFCND1BWP12TLVT (D, E, CP, CDN, Q, QN);
    input D, E, CP, CDN;  
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire D_d, E_d, CP_d ;
    pullup   (SDN);
    tsmc_mux (DE, Q_buf, D_d, E_d);
    tsmc_dff (Q_buf, DE, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (SDN);
    buf      (CDN_i, CDN);
    tsmc_mux (DE, Q_buf, D, E);
    tsmc_dff (Q_buf, DE, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    and  (D_check, CDN_i, E_d);
  `else
    not  (E_int_not, E);
    and  (D_check, CDN_i, E);
  `endif
  and  (CP_check, CDN_i, D_check);
  buf  (E_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFCND2BWP12TLVT (D, E, CP, CDN, Q, QN);
    input D, E, CP, CDN;  
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire D_d, E_d, CP_d ;
    pullup   (SDN);
    tsmc_mux (DE, Q_buf, D_d, E_d);
    tsmc_dff (Q_buf, DE, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (SDN);
    buf      (CDN_i, CDN);
    tsmc_mux (DE, Q_buf, D, E);
    tsmc_dff (Q_buf, DE, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    and  (D_check, CDN_i, E_d);
  `else
    not  (E_int_not, E);
    and  (D_check, CDN_i, E);
  `endif
  and  (CP_check, CDN_i, D_check);
  buf  (E_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFCND4BWP12TLVT (D, E, CP, CDN, Q, QN);
    input D, E, CP, CDN;  
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire D_d, E_d, CP_d ;
    pullup   (SDN);
    tsmc_mux (DE, Q_buf, D_d, E_d);
    tsmc_dff (Q_buf, DE, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (SDN);
    buf      (CDN_i, CDN);
    tsmc_mux (DE, Q_buf, D, E);
    tsmc_dff (Q_buf, DE, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    and  (D_check, CDN_i, E_d);
  `else
    not  (E_int_not, E);
    and  (D_check, CDN_i, E);
  `endif
  and  (CP_check, CDN_i, D_check);
  buf  (E_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFCNQD1BWP12TLVT (D, E, CP, CDN, Q);
    input D, E, CP, CDN;  
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire D_d, E_d, CP_d ;
    pullup   (SDN);
    tsmc_mux (DE, Q_buf, D_d, E_d);
    tsmc_dff (Q_buf, DE, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (SDN);
    buf      (CDN_i, CDN);
    tsmc_mux (DE, Q_buf, D, E);
    tsmc_dff (Q_buf, DE, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    and  (D_check, CDN_i, E_d);
  `else
    not  (E_int_not, E);
    and  (D_check, CDN_i, E);
  `endif
  and  (CP_check, CDN_i, D_check);
  buf  (E_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFCNQD2BWP12TLVT (D, E, CP, CDN, Q);
    input D, E, CP, CDN;  
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire D_d, E_d, CP_d ;
    pullup   (SDN);
    tsmc_mux (DE, Q_buf, D_d, E_d);
    tsmc_dff (Q_buf, DE, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (SDN);
    buf      (CDN_i, CDN);
    tsmc_mux (DE, Q_buf, D, E);
    tsmc_dff (Q_buf, DE, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    and  (D_check, CDN_i, E_d);
  `else
    not  (E_int_not, E);
    and  (D_check, CDN_i, E);
  `endif
  and  (CP_check, CDN_i, D_check);
  buf  (E_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFCNQD4BWP12TLVT (D, E, CP, CDN, Q);
    input D, E, CP, CDN;  
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire D_d, E_d, CP_d ;
    pullup   (SDN);
    tsmc_mux (DE, Q_buf, D_d, E_d);
    tsmc_dff (Q_buf, DE, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (SDN);
    buf      (CDN_i, CDN);
    tsmc_mux (DE, Q_buf, D, E);
    tsmc_dff (Q_buf, DE, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    and  (D_check, CDN_i, E_d);
  `else
    not  (E_int_not, E);
    and  (D_check, CDN_i, E);
  `endif
  and  (CP_check, CDN_i, D_check);
  buf  (E_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFD1BWP12TLVT (D, E, CP, Q, QN);
    input D, E, CP;  
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, E_d, CP_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (DE, Q_buf, D_d, E_d);
    tsmc_dff (Q_buf, DE, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (DE, Q_buf, D, E);
    tsmc_dff (Q_buf, DE, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    buf  (D_check, E_d);
  `else
    not  (E_int_not, E);
    buf  (D_check, E);
  `endif
  buf  (CP_check, D_check);
  pullup  (E_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFD2BWP12TLVT (D, E, CP, Q, QN);
    input D, E, CP;  
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, E_d, CP_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (DE, Q_buf, D_d, E_d);
    tsmc_dff (Q_buf, DE, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (DE, Q_buf, D, E);
    tsmc_dff (Q_buf, DE, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    buf  (D_check, E_d);
  `else
    not  (E_int_not, E);
    buf  (D_check, E);
  `endif
  buf  (CP_check, D_check);
  pullup  (E_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFD4BWP12TLVT (D, E, CP, Q, QN);
    input D, E, CP;  
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, E_d, CP_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (DE, Q_buf, D_d, E_d);
    tsmc_dff (Q_buf, DE, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (DE, Q_buf, D, E);
    tsmc_dff (Q_buf, DE, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    buf  (D_check, E_d);
  `else
    not  (E_int_not, E);
    buf  (D_check, E);
  `endif
  buf  (CP_check, D_check);
  pullup  (E_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFKCND1BWP12TLVT (D, E, CP, CN, Q, QN);
    input D, E, CP, CN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, E_d, CP_d, CN_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    and      (D2, CN_d, D1);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    and      (D2, CN, D1);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (CN_int_not, CN_d);
    buf  (E_check, CN_d);
    and  (D_check, CN_d, E_d);
  `else
    not  (CN_int_not, CN);
    buf  (E_check, CN);
    and  (D_check, CN, E);
  `endif
  or   (CP_check, CN_int_not, D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && E && D) || (CN && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((CN && E && D) || (CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFKCND2BWP12TLVT (D, E, CP, CN, Q, QN);
    input D, E, CP, CN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, E_d, CP_d, CN_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    and      (D2, CN_d, D1);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    and      (D2, CN, D1);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (CN_int_not, CN_d);
    buf  (E_check, CN_d);
    and  (D_check, CN_d, E_d);
  `else
    not  (CN_int_not, CN);
    buf  (E_check, CN);
    and  (D_check, CN, E);
  `endif
  or   (CP_check, CN_int_not, D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && E && D) || (CN && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((CN && E && D) || (CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFKCND4BWP12TLVT (D, E, CP, CN, Q, QN);
    input D, E, CP, CN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, E_d, CP_d, CN_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    and      (D2, CN_d, D1);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    and      (D2, CN, D1);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (CN_int_not, CN_d);
    buf  (E_check, CN_d);
    and  (D_check, CN_d, E_d);
  `else
    not  (CN_int_not, CN);
    buf  (E_check, CN);
    and  (D_check, CN, E);
  `endif
  or   (CP_check, CN_int_not, D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && E && D) || (CN && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((CN && E && D) || (CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFKCNQD1BWP12TLVT (D, E, CP, CN, Q);
    input D, E, CP, CN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, E_d, CP_d, CN_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    and      (D2, CN_d, D1);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    and      (D2, CN, D1);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (CN_int_not, CN_d);
    buf  (E_check, CN_d);
    and  (D_check, CN_d, E_d);
  `else
    not  (CN_int_not, CN);
    buf  (E_check, CN);
    and  (D_check, CN, E);
  `endif
  or   (CP_check, CN_int_not, D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && E && D) || (CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFKCNQD2BWP12TLVT (D, E, CP, CN, Q);
    input D, E, CP, CN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, E_d, CP_d, CN_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    and      (D2, CN_d, D1);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    and      (D2, CN, D1);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (CN_int_not, CN_d);
    buf  (E_check, CN_d);
    and  (D_check, CN_d, E_d);
  `else
    not  (CN_int_not, CN);
    buf  (E_check, CN);
    and  (D_check, CN, E);
  `endif
  or   (CP_check, CN_int_not, D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && E && D) || (CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFKCNQD4BWP12TLVT (D, E, CP, CN, Q);
    input D, E, CP, CN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, E_d, CP_d, CN_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    and      (D2, CN_d, D1);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    and      (D2, CN, D1);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (CN_int_not, CN_d);
    buf  (E_check, CN_d);
    and  (D_check, CN_d, E_d);
  `else
    not  (CN_int_not, CN);
    buf  (E_check, CN);
    and  (D_check, CN, E);
  `endif
  or   (CP_check, CN_int_not, D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((CN && E && D) || (CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFQD1BWP12TLVT (D, E, CP, Q);
    input D, E, CP;  
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, E_d, CP_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (DE, Q_buf, D_d, E_d);
    tsmc_dff (Q_buf, DE, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (DE, Q_buf, D, E);
    tsmc_dff (Q_buf, DE, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    buf  (D_check, E_d);
  `else
    not  (E_int_not, E);
    buf  (D_check, E);
  `endif
  buf  (CP_check, D_check);
  pullup  (E_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFQD2BWP12TLVT (D, E, CP, Q);
    input D, E, CP;  
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, E_d, CP_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (DE, Q_buf, D_d, E_d);
    tsmc_dff (Q_buf, DE, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (DE, Q_buf, D, E);
    tsmc_dff (Q_buf, DE, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    buf  (D_check, E_d);
  `else
    not  (E_int_not, E);
    buf  (D_check, E);
  `endif
  buf  (CP_check, D_check);
  pullup  (E_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module EDFQD4BWP12TLVT (D, E, CP, Q);
    input D, E, CP;  
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, E_d, CP_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (DE, Q_buf, D_d, E_d);
    tsmc_dff (Q_buf, DE, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (DE, Q_buf, D, E);
    tsmc_dff (Q_buf, DE, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    buf  (D_check, E_d);
  `else
    not  (E_int_not, E);
    buf  (D_check, E);
  `endif
  buf  (CP_check, D_check);
  pullup  (E_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((E && D) || (!(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module FA1D0BWP12TLVT (A, B, CI, S, CO);
  input		A, B, CI;
  output	S, CO;
  xor		(S, A, B, CI);
  and		(n2, A, B);
  and		(n3, A, CI);
  and		(n4, B, CI);
  or		(CO, n2, n3, n4);

  specify
    if (B == 1'b0 && CI == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => CO) = (0, 0);
    ifnone (A => CO) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CO) = (0, 0);
    ifnone (B => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CO) = (0, 0);
    ifnone (CI => CO) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    ifnone (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FA1D1BWP12TLVT (A, B, CI, S, CO);
  input		A, B, CI;
  output	S, CO;
  xor		(S, A, B, CI);
  and		(n2, A, B);
  and		(n3, A, CI);
  and		(n4, B, CI);
  or		(CO, n2, n3, n4);

  specify
    if (B == 1'b0 && CI == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => CO) = (0, 0);
    ifnone (A => CO) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CO) = (0, 0);
    ifnone (B => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CO) = (0, 0);
    ifnone (CI => CO) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    ifnone (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FA1D2BWP12TLVT (A, B, CI, S, CO);
  input		A, B, CI;
  output	S, CO;
  xor		(S, A, B, CI);
  and		(n2, A, B);
  and		(n3, A, CI);
  and		(n4, B, CI);
  or		(CO, n2, n3, n4);

  specify
    if (B == 1'b0 && CI == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => CO) = (0, 0);
    ifnone (A => CO) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CO) = (0, 0);
    ifnone (B => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CO) = (0, 0);
    ifnone (CI => CO) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    ifnone (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FA1D4BWP12TLVT (A, B, CI, S, CO);
  input		A, B, CI;
  output	S, CO;
  xor		(S, A, B, CI);
  and		(n2, A, B);
  and		(n3, A, CI);
  and		(n4, B, CI);
  or		(CO, n2, n3, n4);

  specify
    if (B == 1'b0 && CI == 1'b1)
    (A => CO) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => CO) = (0, 0);
    ifnone (A => CO) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CO) = (0, 0);
    ifnone (B => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CO) = (0, 0);
    ifnone (CI => CO) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    ifnone (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FCICIND1BWP12TLVT (A, B, CIN, CO);
input A, B, CIN;
output CO;
  and  (temp1, A, B);
  not  (CINB, CIN);
  and  (temp2, A, CINB);
  and  (temp3, B, CINB);
  or   (CO, temp1, temp2, temp3);

  specify
    if (B == 1'b0 && CIN == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b1 && CIN == 1'b1)
    (A => CO) = (0, 0);
    ifnone (A => CO) = (0, 0);
    if (A == 1'b0 && CIN == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b1 && CIN == 1'b1)
    (B => CO) = (0, 0);
    ifnone (B => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CIN => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CIN => CO) = (0, 0);
    ifnone (CIN => CO) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FCICIND2BWP12TLVT (A, B, CIN, CO);
input A, B, CIN;
output CO;
  and  (temp1, A, B);
  not  (CINB, CIN);
  and  (temp2, A, CINB);
  and  (temp3, B, CINB);
  or   (CO, temp1, temp2, temp3);

  specify
    if (B == 1'b0 && CIN == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b1 && CIN == 1'b1)
    (A => CO) = (0, 0);
    ifnone (A => CO) = (0, 0);
    if (A == 1'b0 && CIN == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b1 && CIN == 1'b1)
    (B => CO) = (0, 0);
    ifnone (B => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CIN => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CIN => CO) = (0, 0);
    ifnone (CIN => CO) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FCICOND1BWP12TLVT (A, B, CI, CON);
input A, B, CI;
output CON;
  and  (temp1, A, B);
  and  (temp2, A, CI);
  and  (temp3, B, CI);
  or   (CO, temp1, temp2, temp3);
  not  (CON, CO);

  specify
    if (B == 1'b0 && CI == 1'b1)
    (A => CON) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => CON) = (0, 0);
    ifnone (A => CON) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CON) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CON) = (0, 0);
    ifnone (B => CON) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CON) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CON) = (0, 0);
    ifnone (CI => CON) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FCICOND2BWP12TLVT (A, B, CI, CON);
input A, B, CI;
output CON;
  and  (temp1, A, B);
  and  (temp2, A, CI);
  and  (temp3, B, CI);
  or   (CO, temp1, temp2, temp3);
  not  (CON, CO);

  specify
    if (B == 1'b0 && CI == 1'b1)
    (A => CON) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => CON) = (0, 0);
    ifnone (A => CON) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CON) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CON) = (0, 0);
    ifnone (B => CON) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CON) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CON) = (0, 0);
    ifnone (CI => CON) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FCSICIND1BWP12TLVT (A, B, CIN0, CIN1, CS, S, CO0, CO1);
   input A, B, CIN0, CIN1, CS;
   output S;
   output CO0 ;
   output CO1 ;
   tsmc_mux (I0_out, CIN0, CIN1, CS);
   xor (I1_out, I0_out, A);
   xor (I2_out, I1_out, B);
   not (S, I2_out);
   not (I4_out, B);
   not (I5_out, A);
   and (I6_out, I4_out, I5_out);
   not (I7_out, A);
   and (I8_out, I7_out, CIN0);
   not (I10_out, B);
   and (I11_out, CIN0, I10_out);
   or  (I12_out, I6_out, I8_out, I11_out);
   not (CO0, I12_out);
   not (I14_out, B);
   not (I15_out, A);
   and (I16_out, I14_out, I15_out);
   not (I17_out, A);
   and (I18_out, I17_out, CIN1);
   not (I20_out, B);
   and (I21_out, CIN1, I20_out);
   or  (I22_out, I16_out, I18_out, I21_out);
   not (CO1, I22_out);

  specify
    if (B == 1'b0 && CIN0 == 1'b0)
    (A => CO0) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1)
    (A => CO0) = (0, 0);
    ifnone (A => CO0) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0)
    (B => CO0) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1)
    (B => CO0) = (0, 0);
    ifnone (B => CO0) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CIN0 => CO0) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CIN0 => CO0) = (0, 0);
    ifnone (CIN0 => CO0) = (0, 0);
    if (B == 1'b0 && CIN1 == 1'b0)
    (A => CO1) = (0, 0);
    if (B == 1'b1 && CIN1 == 1'b1)
    (A => CO1) = (0, 0);
    ifnone (A => CO1) = (0, 0);
    if (A == 1'b0 && CIN1 == 1'b0)
    (B => CO1) = (0, 0);
    if (A == 1'b1 && CIN1 == 1'b1)
    (B => CO1) = (0, 0);
    ifnone (B => CO1) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CIN1 => CO1) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CIN1 => CO1) = (0, 0);
    ifnone (CIN1 => CO1) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    ifnone (CIN0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b0 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b1 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b0 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b1 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN0 == 1'b0 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN0 == 1'b1 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    ifnone (CIN1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1)
    (CS => S) = (0, 0);
    ifnone (CS => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FCSICIND2BWP12TLVT (A, B, CIN0, CIN1, CS, S, CO0, CO1);
   input A, B, CIN0, CIN1, CS;
   output S;
   output CO0 ;
   output CO1 ;
   tsmc_mux (I0_out, CIN0, CIN1, CS);
   xor (I1_out, I0_out, A);
   xor (I2_out, I1_out, B);
   not (S, I2_out);
   not (I4_out, B);
   not (I5_out, A);
   and (I6_out, I4_out, I5_out);
   not (I7_out, A);
   and (I8_out, I7_out, CIN0);
   not (I10_out, B);
   and (I11_out, CIN0, I10_out);
   or  (I12_out, I6_out, I8_out, I11_out);
   not (CO0, I12_out);
   not (I14_out, B);
   not (I15_out, A);
   and (I16_out, I14_out, I15_out);
   not (I17_out, A);
   and (I18_out, I17_out, CIN1);
   not (I20_out, B);
   and (I21_out, CIN1, I20_out);
   or  (I22_out, I16_out, I18_out, I21_out);
   not (CO1, I22_out);

  specify
    if (B == 1'b0 && CIN0 == 1'b0)
    (A => CO0) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1)
    (A => CO0) = (0, 0);
    ifnone (A => CO0) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0)
    (B => CO0) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1)
    (B => CO0) = (0, 0);
    ifnone (B => CO0) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CIN0 => CO0) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CIN0 => CO0) = (0, 0);
    ifnone (CIN0 => CO0) = (0, 0);
    if (B == 1'b0 && CIN1 == 1'b0)
    (A => CO1) = (0, 0);
    if (B == 1'b1 && CIN1 == 1'b1)
    (A => CO1) = (0, 0);
    ifnone (A => CO1) = (0, 0);
    if (A == 1'b0 && CIN1 == 1'b0)
    (B => CO1) = (0, 0);
    if (A == 1'b1 && CIN1 == 1'b1)
    (B => CO1) = (0, 0);
    ifnone (B => CO1) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CIN1 => CO1) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CIN1 => CO1) = (0, 0);
    ifnone (CIN1 => CO1) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN1 == 1'b0 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN1 == 1'b1 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN1 == 1'b0 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN1 == 1'b1 && CS == 1'b0)
    (CIN0 => S) = (0, 0);
    ifnone (CIN0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b0 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CIN0 == 1'b1 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b0 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CIN0 == 1'b1 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN0 == 1'b0 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN0 == 1'b1 && CS == 1'b1)
    (CIN1 => S) = (0, 0);
    ifnone (CIN1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN0 == 1'b1 && CIN1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN0 == 1'b1 && CIN1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CIN0 == 1'b0 && CIN1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CIN0 == 1'b0 && CIN1 == 1'b1)
    (CS => S) = (0, 0);
    ifnone (CS => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FCSICOND1BWP12TLVT (A, B, CI0, CI1, CS, S, CON0, CON1);
   input A, B, CI0, CI1, CS;
   output S;
   output CON0 ;
   output CON1 ;
   tsmc_mux (I0_out, CI0, CI1, CS);
   xor (I1_out, I0_out, A);
   xor (S, I1_out, B);
   and (I3_out, A, B);
   and (I4_out, B, CI0);
   and (I6_out, CI0, A);
   or  (I7_out, I3_out, I4_out, I6_out);
   not (CON0, I7_out);
   and (I9_out, A, B);
   and (I10_out, B, CI1);
   and (I12_out, CI1, A);
   or  (I13_out, I9_out, I10_out, I12_out);
   not (CON1, I13_out);

  specify
    if (B == 1'b0 && CI0 == 1'b1)
    (A => CON0) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0)
    (A => CON0) = (0, 0);
    ifnone (A => CON0) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1)
    (B => CON0) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0)
    (B => CON0) = (0, 0);
    ifnone (B => CON0) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI0 => CON0) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI0 => CON0) = (0, 0);
    ifnone (CI0 => CON0) = (0, 0);
    if (B == 1'b0 && CI1 == 1'b1)
    (A => CON1) = (0, 0);
    if (B == 1'b1 && CI1 == 1'b0)
    (A => CON1) = (0, 0);
    ifnone (A => CON1) = (0, 0);
    if (A == 1'b0 && CI1 == 1'b1)
    (B => CON1) = (0, 0);
    if (A == 1'b1 && CI1 == 1'b0)
    (B => CON1) = (0, 0);
    ifnone (B => CON1) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI1 => CON1) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI1 => CON1) = (0, 0);
    ifnone (CI1 => CON1) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    ifnone (CI0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI0 == 1'b0 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI0 == 1'b1 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b0 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b1 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b0 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b1 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    ifnone (CI1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0)
    (CS => S) = (0, 0);
    ifnone (CS => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FCSICOND2BWP12TLVT (A, B, CI0, CI1, CS, S, CON0, CON1);
   input A, B, CI0, CI1, CS;
   output S;
   output CON0 ;
   output CON1 ;
   tsmc_mux (I0_out, CI0, CI1, CS);
   xor (I1_out, I0_out, A);
   xor (S, I1_out, B);
   and (I3_out, A, B);
   and (I4_out, B, CI0);
   and (I6_out, CI0, A);
   or  (I7_out, I3_out, I4_out, I6_out);
   not (CON0, I7_out);
   and (I9_out, A, B);
   and (I10_out, B, CI1);
   and (I12_out, CI1, A);
   or  (I13_out, I9_out, I10_out, I12_out);
   not (CON1, I13_out);

  specify
    if (B == 1'b0 && CI0 == 1'b1)
    (A => CON0) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0)
    (A => CON0) = (0, 0);
    ifnone (A => CON0) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1)
    (B => CON0) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0)
    (B => CON0) = (0, 0);
    ifnone (B => CON0) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI0 => CON0) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI0 => CON0) = (0, 0);
    ifnone (CI0 => CON0) = (0, 0);
    if (B == 1'b0 && CI1 == 1'b1)
    (A => CON1) = (0, 0);
    if (B == 1'b1 && CI1 == 1'b0)
    (A => CON1) = (0, 0);
    ifnone (A => CON1) = (0, 0);
    if (A == 1'b0 && CI1 == 1'b1)
    (B => CON1) = (0, 0);
    if (A == 1'b1 && CI1 == 1'b0)
    (B => CON1) = (0, 0);
    ifnone (B => CON1) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI1 => CON1) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI1 => CON1) = (0, 0);
    ifnone (CI1 => CON1) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI0 == 1'b1 && CI1 == 1'b1 && CS == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0 && CS == 1'b1)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI1 == 1'b0 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI1 == 1'b1 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI1 == 1'b0 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI1 == 1'b1 && CS == 1'b0)
    (CI0 => S) = (0, 0);
    ifnone (CI0 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI0 == 1'b0 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI0 == 1'b1 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b0 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1 && CI0 == 1'b1 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b0 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0 && CI0 == 1'b1 && CS == 1'b1)
    (CI1 => S) = (0, 0);
    ifnone (CI1 => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI0 == 1'b0 && CI1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI0 == 1'b0 && CI1 == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0 && CI0 == 1'b1 && CI1 == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1 && CI0 == 1'b1 && CI1 == 1'b0)
    (CS => S) = (0, 0);
    ifnone (CS => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FICIND1BWP12TLVT (A, B, CIN, S, CO);
input A, B, CIN;
output S, CO;
  not  (CINB, CIN);
  xor  (S, A, B, CINB);
  and  (temp1, A, B);
  and  (temp2, A, CINB);
  and  (temp3, B, CINB);
  or   (CO, temp1, temp2, temp3);

  specify
    if (B == 1'b0 && CIN == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b1 && CIN == 1'b1)
    (A => CO) = (0, 0);
    ifnone (A => CO) = (0, 0);
    if (A == 1'b0 && CIN == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b1 && CIN == 1'b1)
    (B => CO) = (0, 0);
    ifnone (B => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CIN => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CIN => CO) = (0, 0);
    ifnone (CIN => CO) = (0, 0);
    if (B == 1'b0 && CIN == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN == 1'b1)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0 && CIN == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN == 1'b1)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CIN => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CIN => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CIN => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CIN => S) = (0, 0);
    ifnone (CIN => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FICIND2BWP12TLVT (A, B, CIN, S, CO);
input A, B, CIN;
output S, CO;
  not  (CINB, CIN);
  xor  (S, A, B, CINB);
  and  (temp1, A, B);
  and  (temp2, A, CINB);
  and  (temp3, B, CINB);
  or   (CO, temp1, temp2, temp3);

  specify
    if (B == 1'b0 && CIN == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b1 && CIN == 1'b1)
    (A => CO) = (0, 0);
    ifnone (A => CO) = (0, 0);
    if (A == 1'b0 && CIN == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b1 && CIN == 1'b1)
    (B => CO) = (0, 0);
    ifnone (B => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CIN => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CIN => CO) = (0, 0);
    ifnone (CIN => CO) = (0, 0);
    if (B == 1'b0 && CIN == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CIN == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CIN == 1'b1)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0 && CIN == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CIN == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CIN == 1'b1)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CIN => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CIN => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CIN => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CIN => S) = (0, 0);
    ifnone (CIN => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FICOND1BWP12TLVT (A, B, CI, S, CON);
input A, B, CI;
output S, CON;
  xor  (S, A, B, CI);
  and  (temp1, A, B);
  and  (temp2, A, CI);
  and  (temp3, B, CI);
  or   (CO, temp1, temp2, temp3);
  not  (CON, CO);

  specify
    if (B == 1'b0 && CI == 1'b1)
    (A => CON) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => CON) = (0, 0);
    ifnone (A => CON) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CON) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CON) = (0, 0);
    ifnone (B => CON) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CON) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CON) = (0, 0);
    ifnone (CI => CON) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    ifnone (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FICOND2BWP12TLVT (A, B, CI, S, CON);
input A, B, CI;
output S, CON;
  xor  (S, A, B, CI);
  and  (temp1, A, B);
  and  (temp2, A, CI);
  and  (temp3, B, CI);
  or   (CO, temp1, temp2, temp3);
  not  (CON, CO);

  specify
    if (B == 1'b0 && CI == 1'b1)
    (A => CON) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => CON) = (0, 0);
    ifnone (A => CON) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CON) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CON) = (0, 0);
    ifnone (B => CON) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CON) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CON) = (0, 0);
    ifnone (CI => CON) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    ifnone (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FIICOND1BWP12TLVT (A, B, C, S, CON0, CON1);
input A, B, C;
output S, CON0, CON1;
  xor  (S, A, B, C);
  and  (temp1, A, B);
  or   (temp2, A, B);
  not  (CON0, temp1);
  not  (CON1, temp2);

  specify
    (A => CON0) = (0, 0);
    (B => CON0) = (0, 0);
    (A => CON1) = (0, 0);
    (B => CON1) = (0, 0);
    if (B == 1'b0 && C == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0 && C == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (C => S) = (0, 0);
    ifnone (C => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FIICOND2BWP12TLVT (A, B, C, S, CON0, CON1);
input A, B, C;
output S, CON0, CON1;
  xor  (S, A, B, C);
  and  (temp1, A, B);
  or   (temp2, A, B);
  not  (CON0, temp1);
  not  (CON1, temp2);

  specify
    (A => CON0) = (0, 0);
    (B => CON0) = (0, 0);
    (A => CON1) = (0, 0);
    (B => CON1) = (0, 0);
    if (B == 1'b0 && C == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && C == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b1 && C == 1'b0)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0 && C == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && C == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && C == 1'b0)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (C => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (C => S) = (0, 0);
    ifnone (C => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GAN2D1BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GAN2D2BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GAOI21D1BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and		(A, A1, A2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GAOI21D2BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and		(A, A1, A2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GAOI22D1BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and		(A, A1, A2);
    and		(B, B1, B2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFD1BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFD2BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFD3BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFD4BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFD8BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GDCAP10BWP12TLVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GDCAP2BWP12TLVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GDCAP3BWP12TLVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GDCAP4BWP12TLVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GDCAPBWP12TLVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GDFCNQD1BWP12TLVT (D, CP, CDN, Q);
    input D, CP, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire D_d, CP_d ;
    pullup   (SDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    pullup   (SDN);
    tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (CP_check, CDN_i);
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module GDFQD1BWP12TLVT (D, CP, Q);
    input D, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, CP_d ;
    pullup	 (CDN);
    pullup	 (SDN);
    tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup	 (CDN);
    pullup	 (SDN);
    tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  pullup  (CP_check);
  pullup  (D_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:D)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module GFILL10BWP12TLVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GFILL2BWP12TLVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GFILL3BWP12TLVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GFILL4BWP12TLVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GFILLBWP12TLVT;
    // No function
endmodule
`endcelldefine



`celldefine
module GINVD1BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GINVD2BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GINVD3BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GINVD4BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GINVD8BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GMUX2D1BWP12TLVT (I0, I1, S, Z);
   input S, I1, I0;
   output Z;
   tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    ifnone (I0 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    ifnone (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
    ifnone (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GMUX2D2BWP12TLVT (I0, I1, S, Z);
   input S, I1, I0;
   output Z;
   tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    ifnone (I0 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    ifnone (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
    ifnone (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GMUX2ND1BWP12TLVT (I0, I1, S, ZN);
   input I0, I1, S;
   output ZN;
   tsmc_mux (I0_out, I0, I1, S);
   not (ZN, I0_out);

  specify
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    ifnone (I0 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    ifnone (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
    ifnone (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GMUX2ND2BWP12TLVT (I0, I1, S, ZN);
   input I0, I1, S;
   output ZN;
   tsmc_mux (I0_out, I0, I1, S);
   not (ZN, I0_out);

  specify
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    ifnone (I0 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    ifnone (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
    ifnone (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND2D1BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nand		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND2D2BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nand		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND2D3BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nand		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND2D4BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nand		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND3D1BWP12TLVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    nand		(ZN, A1, A2, A3);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND3D2BWP12TLVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    nand		(ZN, A1, A2, A3);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GNR2D1BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nor		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GNR2D2BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nor		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GNR3D1BWP12TLVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    nor		(ZN, A1, A2, A3);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GNR3D2BWP12TLVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    nor		(ZN, A1, A2, A3);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GOAI21D1BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or		(A, A1, A2);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GOAI21D2BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or		(A, A1, A2);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GOR2D1BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GOR2D2BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GSDFCNQD1BWP12TLVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    pullup       (SDN);
    tsmc_mux     (D_i, D_d, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CP_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module GTIEHBWP12TLVT (Z);
  output  Z;
  buf (Z, 1'b1);

endmodule
`endcelldefine

`celldefine
module GTIELBWP12TLVT (ZN);
  output  ZN;
  buf (ZN, 1'b0);

endmodule
`endcelldefine

`celldefine
module GXNR2D1BWP12TLVT (A1, A2, ZN);
  input		A1, A2;
  output 	ZN;
  xnor		(ZN, A1, A2);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    ifnone (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
    ifnone (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GXNR2D2BWP12TLVT (A1, A2, ZN);
  input		A1, A2;
  output 	ZN;
  xnor		(ZN, A1, A2);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    ifnone (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
    ifnone (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GXOR2D1BWP12TLVT (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
  xor		(Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    ifnone (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
    ifnone (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GXOR2D2BWP12TLVT (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
  xor		(Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    ifnone (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
    ifnone (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HA1D0BWP12TLVT (A, B, S, CO);
  input	 	A, B;
  output	S, CO;
  xor		(S, A, B);
  and		(CO, A, B);

  specify
    (A => CO) = (0, 0);
    (B => CO) = (0, 0);
    if (B == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HA1D1BWP12TLVT (A, B, S, CO);
  input	 	A, B;
  output	S, CO;
  xor		(S, A, B);
  and		(CO, A, B);

  specify
    (A => CO) = (0, 0);
    (B => CO) = (0, 0);
    if (B == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HA1D2BWP12TLVT (A, B, S, CO);
  input	 	A, B;
  output	S, CO;
  xor		(S, A, B);
  and		(CO, A, B);

  specify
    (A => CO) = (0, 0);
    (B => CO) = (0, 0);
    if (B == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HA1D4BWP12TLVT (A, B, S, CO);
  input	 	A, B;
  output	S, CO;
  xor		(S, A, B);
  and		(CO, A, B);

  specify
    (A => CO) = (0, 0);
    (B => CO) = (0, 0);
    if (B == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1)
    (B => S) = (0, 0);
    ifnone (B => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HCOSCIND1BWP12TLVT (A, CIN, CS, S, CO);
   input A, CIN, CS;
   output S;
   output CO ;
   xor (I0_out, A, CIN);
   not (I1_out, I0_out);
   tsmc_mux (S, A, I1_out, CS);
   not (I3_out, CIN);
   and (CO, I3_out, A);

  specify
    (A => CO) = (0, 0);
    (CIN => CO) = (0, 0);
    if (CIN == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (CIN == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (CIN == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (CIN == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b1 && CS == 1'b1)
    (CIN => S) = (0, 0);
    if (A == 1'b0 && CS == 1'b1)
    (CIN => S) = (0, 0);
    ifnone (CIN => S) = (0, 0);
    if (A == 1'b0 && CIN == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b1 && CIN == 1'b0)
    (CS => S) = (0, 0);
    ifnone (CS => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HCOSCIND2BWP12TLVT (A, CIN, CS, S, CO);
   input A, CIN, CS;
   output S;
   output CO ;
   xor (I0_out, A, CIN);
   not (I1_out, I0_out);
   tsmc_mux (S, A, I1_out, CS);
   not (I3_out, CIN);
   and (CO, I3_out, A);

  specify
    (A => CO) = (0, 0);
    (CIN => CO) = (0, 0);
    if (CIN == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (CIN == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (CIN == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    if (CIN == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b1 && CS == 1'b1)
    (CIN => S) = (0, 0);
    if (A == 1'b0 && CS == 1'b1)
    (CIN => S) = (0, 0);
    ifnone (CIN => S) = (0, 0);
    if (A == 1'b0 && CIN == 1'b0)
    (CS => S) = (0, 0);
    if (A == 1'b1 && CIN == 1'b0)
    (CS => S) = (0, 0);
    ifnone (CS => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HCOSCOND1BWP12TLVT (A, CI, CS, S, CON);
   input A, CI, CS;
   output S;
   output CON ;
   xor (I0_out, A, CI);
   tsmc_mux (S, A, I0_out, CS);
   and (I2_out, A, CI);
   not (CON, I2_out);

  specify
    (A => CON) = (0, 0);
    (CI => CON) = (0, 0);
    if (CI == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (CI == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (CI == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (CI == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0 && CS == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b1 && CS == 1'b1)
    (CI => S) = (0, 0);
    ifnone (CI => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (CS => S) = (0, 0);
    ifnone (CS => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HCOSCOND2BWP12TLVT (A, CI, CS, S, CON);
   input A, CI, CS;
   output S;
   output CON ;
   xor (I0_out, A, CI);
   tsmc_mux (S, A, I0_out, CS);
   and (I2_out, A, CI);
   not (CON, I2_out);

  specify
    (A => CON) = (0, 0);
    (CI => CON) = (0, 0);
    if (CI == 1'b0 && CS == 1'b0)
    (A => S) = (0, 0);
    if (CI == 1'b0 && CS == 1'b1)
    (A => S) = (0, 0);
    if (CI == 1'b1 && CS == 1'b0)
    (A => S) = (0, 0);
    if (CI == 1'b1 && CS == 1'b1)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0 && CS == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b1 && CS == 1'b1)
    (CI => S) = (0, 0);
    ifnone (CI => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (CS => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (CS => S) = (0, 0);
    ifnone (CS => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HICIND1BWP12TLVT (A, CIN, S, CO);
input A, CIN;
output S, CO;
  not  (CINB, CIN);
  xor  (S, A, CINB);
  and  (CO, A, CINB);

  specify
    (A => CO) = (0, 0);
    (CIN => CO) = (0, 0);
    if (CIN == 1'b1)
    (A => S) = (0, 0);
    if (CIN == 1'b0)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b1)
    (CIN => S) = (0, 0);
    if (A == 1'b0)
    (CIN => S) = (0, 0);
    ifnone (CIN => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HICIND2BWP12TLVT (A, CIN, S, CO);
input A, CIN;
output S, CO;
  not  (CINB, CIN);
  xor  (S, A, CINB);
  and  (CO, A, CINB);

  specify
    (A => CO) = (0, 0);
    (CIN => CO) = (0, 0);
    if (CIN == 1'b1)
    (A => S) = (0, 0);
    if (CIN == 1'b0)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b1)
    (CIN => S) = (0, 0);
    if (A == 1'b0)
    (CIN => S) = (0, 0);
    ifnone (CIN => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HICOND1BWP12TLVT (A, CI, S, CON);
input A, CI;
output S, CON;
  xor  (S, A, CI);
  and  (CO, A, CI);
  not  (CON, CO);

  specify
    (A => CON) = (0, 0);
    (CI => CON) = (0, 0);
    if (CI == 1'b0)
    (A => S) = (0, 0);
    if (CI == 1'b1)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1)
    (CI => S) = (0, 0);
    ifnone (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HICOND2BWP12TLVT (A, CI, S, CON);
input A, CI;
output S, CON;
  xor  (S, A, CI);
  and  (CO, A, CI);
  not  (CON, CO);

  specify
    (A => CON) = (0, 0);
    (CI => CON) = (0, 0);
    if (CI == 1'b0)
    (A => S) = (0, 0);
    if (CI == 1'b1)
    (A => S) = (0, 0);
    ifnone (A => S) = (0, 0);
    if (A == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1)
    (CI => S) = (0, 0);
    ifnone (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IAO21D0BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    not    	(A1N,A1);
    not         (A2N,A2);
    and		(A,A1N,A2N);
    nor         (ZN,A,B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IAO21D1BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    not    	(A1N,A1);
    not         (A2N,A2);
    and		(A,A1N,A2N);
    nor         (ZN,A,B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IAO21D2BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    not    	(A1N,A1);
    not         (A2N,A2);
    and		(A,A1N,A2N);
    nor         (ZN,A,B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IAO21D4BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    not    	(A1N,A1);
    not         (A2N,A2);
    and		(A,A1N,A2N);
    nor         (ZN,A,B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IAO22D0BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not 	(A1N,A1);
    not         (A2N,A2);
    and		(A,A1N,A2N);
    and		(B,B1,B2);
    nor		(ZN,A,B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IAO22D1BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not 	(A1N,A1);
    not         (A2N,A2);
    and		(A,A1N,A2N);
    and		(B,B1,B2);
    nor		(ZN,A,B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IAO22D2BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not 	(A1N,A1);
    not         (A2N,A2);
    and		(A,A1N,A2N);
    and		(B,B1,B2);
    nor		(ZN,A,B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IAO22D4BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not 	(A1N,A1);
    not         (A2N,A2);
    and		(A,A1N,A2N);
    and		(B,B1,B2);
    nor		(ZN,A,B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IIND4D0BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not		    (A1N, A1);
    not         (A2N, A2);
    nand		(ZN, A1N, A2N, B1, B2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IIND4D1BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not		    (A1N, A1);
    not         (A2N, A2);
    nand		(ZN, A1N, A2N, B1, B2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IIND4D2BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not		    (A1N, A1);
    not         (A2N, A2);
    nand		(ZN, A1N, A2N, B1, B2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IIND4D4BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not		    (A1N, A1);
    not         (A2N, A2);
    nand		(ZN, A1N, A2N, B1, B2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IINR4D0BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not		(A1N, A1);
    not     (A2N, A2);
    nor		(ZN, A1N, A2N, B1, B2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IINR4D1BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not		(A1N, A1);
    not     (A2N, A2);
    nor		(ZN, A1N, A2N, B1, B2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IINR4D2BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not		(A1N, A1);
    not     (A2N, A2);
    nor		(ZN, A1N, A2N, B1, B2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IINR4D4BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not		(A1N, A1);
    not     (A2N, A2);
    nor		(ZN, A1N, A2N, B1, B2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND2D0BWP12TLVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not		(A1N, A1);
    nand		(ZN, A1N, B1);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND2D1BWP12TLVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not		(A1N, A1);
    nand		(ZN, A1N, B1);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND2D2BWP12TLVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not		(A1N, A1);
    nand		(ZN, A1N, B1);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND2D4BWP12TLVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not		(A1N, A1);
    nand		(ZN, A1N, B1);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND3D0BWP12TLVT (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not		(A1N, A1);
    nand		(ZN, A1N, B1, B2);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND3D1BWP12TLVT (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not		(A1N, A1);
    nand		(ZN, A1N, B1, B2);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND3D2BWP12TLVT (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not		(A1N, A1);
    nand		(ZN, A1N, B1, B2);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND3D4BWP12TLVT (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not		(A1N, A1);
    nand		(ZN, A1N, B1, B2);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND4D0BWP12TLVT (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not		    (A1N, A1);
    nand		(ZN, A1N, B1, B2, B3);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND4D1BWP12TLVT (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not		    (A1N, A1);
    nand		(ZN, A1N, B1, B2, B3);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND4D2BWP12TLVT (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not		    (A1N, A1);
    nand		(ZN, A1N, B1, B2, B3);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND4D4BWP12TLVT (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not		    (A1N, A1);
    nand		(ZN, A1N, B1, B2, B3);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2D0BWP12TLVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not		(A1N, A1);
    nor		(ZN, A1N, B1);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2D1BWP12TLVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not		(A1N, A1);
    nor		(ZN, A1N, B1);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2D2BWP12TLVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not		(A1N, A1);
    nor		(ZN, A1N, B1);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2D4BWP12TLVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not		(A1N, A1);
    nor		(ZN, A1N, B1);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2XD0BWP12TLVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not		(A1N, A1);
    nor		(ZN, A1N, B1);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2XD1BWP12TLVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not		(A1N, A1);
    nor		(ZN, A1N, B1);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2XD2BWP12TLVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not		(A1N, A1);
    nor		(ZN, A1N, B1);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2XD4BWP12TLVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not		(A1N, A1);
    nor		(ZN, A1N, B1);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR3D0BWP12TLVT (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not		(A1N, A1);
    nor		(ZN, A1N, B1, B2);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR3D1BWP12TLVT (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not		(A1N, A1);
    nor		(ZN, A1N, B1, B2);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR3D2BWP12TLVT (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not		(A1N, A1);
    nor		(ZN, A1N, B1, B2);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR3D4BWP12TLVT (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not		(A1N, A1);
    nor		(ZN, A1N, B1, B2);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR4D0BWP12TLVT (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not		(A1N, A1);
    nor		(ZN, A1N, B1, B2, B3);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR4D1BWP12TLVT (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not		(A1N, A1);
    nor		(ZN, A1N, B1, B2, B3);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR4D2BWP12TLVT (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not		(A1N, A1);
    nor		(ZN, A1N, B1, B2, B3);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR4D4BWP12TLVT (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not		(A1N, A1);
    nor		(ZN, A1N, B1, B2, B3);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD0BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD12BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD16BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD1BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD20BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD24BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD2BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD3BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD4BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD6BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD8BWP12TLVT (I, ZN);
    input I;
    output ZN;
    not		(ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IOA21D0BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    not          (A1N,A1);
    not          (A2N,A2);
    or           (A,A1N,A2N);
    nand         (ZN,A,B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IOA21D1BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    not          (A1N,A1);
    not          (A2N,A2);
    or           (A,A1N,A2N);
    nand         (ZN,A,B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IOA21D2BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    not          (A1N,A1);
    not          (A2N,A2);
    or           (A,A1N,A2N);
    nand         (ZN,A,B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IOA21D4BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    not          (A1N,A1);
    not          (A2N,A2);
    or           (A,A1N,A2N);
    nand         (ZN,A,B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IOA22D0BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not         (A1N,A1);
    not         (A2N,A2);
    or          (A,A1N,A2N);
    or		(B,B1,B2);
    nand        (ZN,A,B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IOA22D1BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not         (A1N,A1);
    not         (A2N,A2);
    or          (A,A1N,A2N);
    or		(B,B1,B2);
    nand        (ZN,A,B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IOA22D2BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not         (A1N,A1);
    not         (A2N,A2);
    or          (A,A1N,A2N);
    or		(B,B1,B2);
    nand        (ZN,A,B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IOA22D4BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    not         (A1N,A1);
    not         (A2N,A2);
    or          (A,A1N,A2N);
    or		(B,B1,B2);
    nand        (ZN,A,B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LHCND1BWP12TLVT (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, E_d ;
    pullup	(SDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup	(SDN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E, 0, notifier);
      $hold (negedge E, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E, 0, notifier);
    $hold (negedge E, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCND2BWP12TLVT (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, E_d ;
    pullup	(SDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup	(SDN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E, 0, notifier);
      $hold (negedge E, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E, 0, notifier);
    $hold (negedge E, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCND4BWP12TLVT (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, E_d ;
    pullup	(SDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup	(SDN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E, 0, notifier);
      $hold (negedge E, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E, 0, notifier);
    $hold (negedge E, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCNDD1BWP12TLVT (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, E_d ;
    pullup	(SDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup	(SDN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E, 0, notifier);
      $hold (negedge E, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E, 0, notifier);
    $hold (negedge E, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCNDD2BWP12TLVT (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, E_d ;
    pullup	(SDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup	(SDN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E, 0, notifier);
      $hold (negedge E, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E, 0, notifier);
    $hold (negedge E, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCNDD4BWP12TLVT (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, E_d ;
    pullup	(SDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup	(SDN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E, 0, notifier);
      $hold (negedge E, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E, 0, notifier);
    $hold (negedge E, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCNDQD1BWP12TLVT (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, E_d ;
    pullup	(SDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup	(SDN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E, 0, notifier);
      $hold (negedge E, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E, 0, notifier);
    $hold (negedge E, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCNDQD2BWP12TLVT (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, E_d ;
    pullup	(SDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup	(SDN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E, 0, notifier);
      $hold (negedge E, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E, 0, notifier);
    $hold (negedge E, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCNDQD4BWP12TLVT (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, E_d ;
    pullup	(SDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup	(SDN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E, 0, notifier);
      $hold (negedge E, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E, 0, notifier);
    $hold (negedge E, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCNQD1BWP12TLVT (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, E_d ;
    pullup	(SDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup	(SDN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E, 0, notifier);
      $hold (negedge E, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E, 0, notifier);
    $hold (negedge E, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCNQD2BWP12TLVT (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, E_d ;
    pullup	(SDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup	(SDN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E, 0, notifier);
      $hold (negedge E, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E, 0, notifier);
    $hold (negedge E, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCNQD4BWP12TLVT (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, E_d ;
    pullup	(SDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup	(SDN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E, 0, notifier);
      $hold (negedge E, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E, 0, notifier);
    $hold (negedge E, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSND1BWP12TLVT (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not		 (QN_buf, Q_buf);
    and		 (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not		 (QN_buf, Q_buf);
    and		 (QN, QN_buf, SDN_i);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E &&& E_DEFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
      $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
    $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSND2BWP12TLVT (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not		 (QN_buf, Q_buf);
    and		 (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not		 (QN_buf, Q_buf);
    and		 (QN, QN_buf, SDN_i);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E &&& E_DEFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
      $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
    $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSND4BWP12TLVT (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not		 (QN_buf, Q_buf);
    and		 (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not		 (QN_buf, Q_buf);
    and		 (QN, QN_buf, SDN_i);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E &&& E_DEFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
      $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
    $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSNDD1BWP12TLVT (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not		 (QN_buf, Q_buf);
    and		 (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not		 (QN_buf, Q_buf);
    and		 (QN, QN_buf, SDN_i);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E &&& E_DEFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
      $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
    $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSNDD2BWP12TLVT (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not		 (QN_buf, Q_buf);
    and		 (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not		 (QN_buf, Q_buf);
    and		 (QN, QN_buf, SDN_i);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E &&& E_DEFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
      $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
    $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSNDD4BWP12TLVT (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not		 (QN_buf, Q_buf);
    and		 (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not		 (QN_buf, Q_buf);
    and		 (QN, QN_buf, SDN_i);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E &&& E_DEFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
      $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
    $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSNDQD1BWP12TLVT (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E &&& E_DEFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
      $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
    $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSNDQD2BWP12TLVT (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E &&& E_DEFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
      $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
    $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSNDQD4BWP12TLVT (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E &&& E_DEFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
      $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
    $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSNQD1BWP12TLVT (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E &&& E_DEFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
      $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
    $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSNQD2BWP12TLVT (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E &&& E_DEFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
      $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
    $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSNQD4BWP12TLVT (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN, negedge E &&& E_DEFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
      $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, negedge E &&& E_DEFCHK, 0, notifier);
    $hold (negedge E &&& E_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHD1BWP12TLVT (D, E, Q, QN);
    input D, E;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, E_d ;
    pullup	 (CDN);
    pullup	 (SDN);
    tsmc_dla (Q_buf, D_d, E_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup	 (CDN);
    pullup	 (SDN);
    tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `endif



  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (posedge E, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge E, posedge D, 0, 0, notifier,,, E_d, D_d);
    $setuphold (negedge E, negedge D, 0, 0, notifier,,, E_d, D_d);
  `else
    $setuphold (negedge E, posedge D, 0, 0, notifier);
    $setuphold (negedge E, negedge D, 0, 0, notifier);
  `endif
  endspecify
endmodule
`endcelldefine

`celldefine
module LHD2BWP12TLVT (D, E, Q, QN);
    input D, E;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, E_d ;
    pullup	 (CDN);
    pullup	 (SDN);
    tsmc_dla (Q_buf, D_d, E_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup	 (CDN);
    pullup	 (SDN);
    tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `endif



  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (posedge E, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge E, posedge D, 0, 0, notifier,,, E_d, D_d);
    $setuphold (negedge E, negedge D, 0, 0, notifier,,, E_d, D_d);
  `else
    $setuphold (negedge E, posedge D, 0, 0, notifier);
    $setuphold (negedge E, negedge D, 0, 0, notifier);
  `endif
  endspecify
endmodule
`endcelldefine

`celldefine
module LHD4BWP12TLVT (D, E, Q, QN);
    input D, E;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, E_d ;
    pullup	 (CDN);
    pullup	 (SDN);
    tsmc_dla (Q_buf, D_d, E_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup	 (CDN);
    pullup	 (SDN);
    tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `endif



  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (posedge E, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge E, posedge D, 0, 0, notifier,,, E_d, D_d);
    $setuphold (negedge E, negedge D, 0, 0, notifier,,, E_d, D_d);
  `else
    $setuphold (negedge E, posedge D, 0, 0, notifier);
    $setuphold (negedge E, negedge D, 0, 0, notifier);
  `endif
  endspecify
endmodule
`endcelldefine

`celldefine
module LHQD1BWP12TLVT (D, E, Q);
    input D, E;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, E_d ;
    pullup	(CDN);
    pullup	(SDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup	(CDN);
    pullup	(SDN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (posedge E, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge E, posedge D, 0, 0, notifier,,, E_d, D_d);
    $setuphold (negedge E, negedge D, 0, 0, notifier,,, E_d, D_d);
  `else
    $setuphold (negedge E, posedge D, 0, 0, notifier);
    $setuphold (negedge E, negedge D, 0, 0, notifier);
  `endif
  endspecify
endmodule
`endcelldefine

`celldefine
module LHQD2BWP12TLVT (D, E, Q);
    input D, E;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, E_d ;
    pullup	(CDN);
    pullup	(SDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup	(CDN);
    pullup	(SDN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (posedge E, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge E, posedge D, 0, 0, notifier,,, E_d, D_d);
    $setuphold (negedge E, negedge D, 0, 0, notifier,,, E_d, D_d);
  `else
    $setuphold (negedge E, posedge D, 0, 0, notifier);
    $setuphold (negedge E, negedge D, 0, 0, notifier);
  `endif
  endspecify
endmodule
`endcelldefine

`celldefine
module LHQD4BWP12TLVT (D, E, Q);
    input D, E;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, E_d ;
    pullup	(CDN);
    pullup	(SDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup	(CDN);
    pullup	(SDN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (posedge E, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge E, posedge D, 0, 0, notifier,,, E_d, D_d);
    $setuphold (negedge E, negedge D, 0, 0, notifier,,, E_d, D_d);
  `else
    $setuphold (negedge E, posedge D, 0, 0, notifier);
    $setuphold (negedge E, negedge D, 0, 0, notifier);
  `endif
  endspecify
endmodule
`endcelldefine

`celldefine
module LHSND1BWP12TLVT (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    pullup	(CDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
    not		(QN_buf, Q_buf);
    and		(QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup	(CDN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
    not		(QN_buf, Q_buf);
    and		(QN, QN_buf, SDN_i);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSND2BWP12TLVT (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    pullup	(CDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
    not		(QN_buf, Q_buf);
    and		(QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup	(CDN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
    not		(QN_buf, Q_buf);
    and		(QN, QN_buf, SDN_i);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSND4BWP12TLVT (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    pullup	(CDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
    not		(QN_buf, Q_buf);
    and		(QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup	(CDN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
    not		(QN_buf, Q_buf);
    and		(QN, QN_buf, SDN_i);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSNDD1BWP12TLVT (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    pullup	(CDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
    not		(QN_buf, Q_buf);
    and		(QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup	(CDN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
    not		(QN_buf, Q_buf);
    and		(QN, QN_buf, SDN_i);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSNDD2BWP12TLVT (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    pullup	(CDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
    not		(QN_buf, Q_buf);
    and		(QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup	(CDN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
    not		(QN_buf, Q_buf);
    and		(QN, QN_buf, SDN_i);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSNDD4BWP12TLVT (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    pullup	(CDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
    not		(QN_buf, Q_buf);
    and		(QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup	(CDN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
    not		(QN_buf, Q_buf);
    and		(QN, QN_buf, SDN_i);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSNDQD1BWP12TLVT (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    pullup	(CDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup	(CDN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSNDQD2BWP12TLVT (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    pullup	(CDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup	(CDN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSNDQD4BWP12TLVT (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    pullup	(CDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup	(CDN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSNQD1BWP12TLVT (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    pullup	(CDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup	(CDN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSNQD2BWP12TLVT (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    pullup	(CDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup	(CDN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSNQD4BWP12TLVT (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, E_d ;
    pullup	(CDN);
    tsmc_dla	(Q_buf, D_d, E_d, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup	(CDN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf         (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (E_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (posedge E, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN, negedge E, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN, negedge E, 0, notifier);
      $hold (negedge E, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge E &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, negedge E, 0, notifier);
    $hold (negedge E, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCND1BWP12TLVT (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, EN_d ;
    pullup       (SDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup       (SDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCND2BWP12TLVT (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, EN_d ;
    pullup       (SDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup       (SDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCND4BWP12TLVT (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, EN_d ;
    pullup       (SDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup       (SDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCNDD1BWP12TLVT (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, EN_d ;
    pullup       (SDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup       (SDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCNDD2BWP12TLVT (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, EN_d ;
    pullup       (SDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup       (SDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCNDD4BWP12TLVT (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, EN_d ;
    pullup       (SDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup       (SDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCNDQD1BWP12TLVT (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, EN_d ;
    pullup       (SDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup       (SDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCNDQD2BWP12TLVT (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, EN_d ;
    pullup       (SDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup       (SDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCNDQD4BWP12TLVT (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, EN_d ;
    pullup       (SDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup       (SDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCNQD1BWP12TLVT (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, EN_d ;
    pullup       (SDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup       (SDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCNQD2BWP12TLVT (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, EN_d ;
    pullup       (SDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup       (SDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCNQD4BWP12TLVT (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire D_d, EN_d ;
    pullup       (SDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup       (SDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSND1BWP12TLVT (D, EN, CDN, SDN, Q, QN);
   input D, EN, CDN, SDN;
   output Q, QN;
   reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
     buf      (CDN_i, CDN_d);
     buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
     buf      (CDN_i, CDN);
     buf      (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
   not		(E, EN_d);
   tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN_i, notifier);
   buf      (Q, Q_buf);
   not		(QN_buf, Q_buf);
   and		(QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
   buf      (CDN_i, CDN);
   buf      (SDN_i, SDN);
   not		(E, EN);
   tsmc_dla	(Q_buf, D, E, CDN_i, SDN_i, notifier);
   buf      (Q, Q_buf);
   not		(QN_buf, Q_buf);
   and		(QN, QN_buf, SDN_i);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN &&& EN_DEFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
      $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
    $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSND2BWP12TLVT (D, EN, CDN, SDN, Q, QN);
   input D, EN, CDN, SDN;
   output Q, QN;
   reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
     buf      (CDN_i, CDN_d);
     buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
     buf      (CDN_i, CDN);
     buf      (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
   not		(E, EN_d);
   tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN_i, notifier);
   buf      (Q, Q_buf);
   not		(QN_buf, Q_buf);
   and		(QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
   buf      (CDN_i, CDN);
   buf      (SDN_i, SDN);
   not		(E, EN);
   tsmc_dla	(Q_buf, D, E, CDN_i, SDN_i, notifier);
   buf      (Q, Q_buf);
   not		(QN_buf, Q_buf);
   and		(QN, QN_buf, SDN_i);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN &&& EN_DEFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
      $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
    $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSND4BWP12TLVT (D, EN, CDN, SDN, Q, QN);
   input D, EN, CDN, SDN;
   output Q, QN;
   reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
     buf      (CDN_i, CDN_d);
     buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
     buf      (CDN_i, CDN);
     buf      (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
   not		(E, EN_d);
   tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN_i, notifier);
   buf      (Q, Q_buf);
   not		(QN_buf, Q_buf);
   and		(QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
   buf      (CDN_i, CDN);
   buf      (SDN_i, SDN);
   not		(E, EN);
   tsmc_dla	(Q_buf, D, E, CDN_i, SDN_i, notifier);
   buf      (Q, Q_buf);
   not		(QN_buf, Q_buf);
   and		(QN, QN_buf, SDN_i);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN &&& EN_DEFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
      $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
    $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSNDD1BWP12TLVT (D, EN, CDN, SDN, Q, QN);
   input D, EN, CDN, SDN;
   output Q, QN;
   reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
     buf      (CDN_i, CDN_d);
     buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
     buf      (CDN_i, CDN);
     buf      (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
   not		(E, EN_d);
   tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN_i, notifier);
   buf      (Q, Q_buf);
   not		(QN_buf, Q_buf);
   and		(QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
   buf      (CDN_i, CDN);
   buf      (SDN_i, SDN);
   not		(E, EN);
   tsmc_dla	(Q_buf, D, E, CDN_i, SDN_i, notifier);
   buf      (Q, Q_buf);
   not		(QN_buf, Q_buf);
   and		(QN, QN_buf, SDN_i);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN &&& EN_DEFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
      $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
    $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSNDD2BWP12TLVT (D, EN, CDN, SDN, Q, QN);
   input D, EN, CDN, SDN;
   output Q, QN;
   reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
     buf      (CDN_i, CDN_d);
     buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
     buf      (CDN_i, CDN);
     buf      (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
   not		(E, EN_d);
   tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN_i, notifier);
   buf      (Q, Q_buf);
   not		(QN_buf, Q_buf);
   and		(QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
   buf      (CDN_i, CDN);
   buf      (SDN_i, SDN);
   not		(E, EN);
   tsmc_dla	(Q_buf, D, E, CDN_i, SDN_i, notifier);
   buf      (Q, Q_buf);
   not		(QN_buf, Q_buf);
   and		(QN, QN_buf, SDN_i);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN &&& EN_DEFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
      $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
    $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSNDD4BWP12TLVT (D, EN, CDN, SDN, Q, QN);
   input D, EN, CDN, SDN;
   output Q, QN;
   reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
     buf      (CDN_i, CDN_d);
     buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
     buf      (CDN_i, CDN);
     buf      (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
   not		(E, EN_d);
   tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN_i, notifier);
   buf      (Q, Q_buf);
   not		(QN_buf, Q_buf);
   and		(QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
   buf      (CDN_i, CDN);
   buf      (SDN_i, SDN);
   not		(E, EN);
   tsmc_dla	(Q_buf, D, E, CDN_i, SDN_i, notifier);
   buf      (Q, Q_buf);
   not		(QN_buf, Q_buf);
   and		(QN, QN_buf, SDN_i);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (CDN => QN) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN &&& EN_DEFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
      $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
    $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSNDQD1BWP12TLVT (D, EN, CDN, SDN, Q);
   input D, EN, CDN, SDN;
   output Q;
   reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
     buf      (CDN_i, CDN_d);
     buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
     buf      (CDN_i, CDN);
     buf      (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
   not		(E, EN_d);
   tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN_i, notifier);
   buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
   buf      (CDN_i, CDN);
   buf      (SDN_i, SDN);
   not		(E, EN);
   tsmc_dla	(Q_buf, D, E, CDN_i, SDN_i, notifier);
   buf          (Q, Q_buf);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN &&& EN_DEFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
      $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
    $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSNDQD2BWP12TLVT (D, EN, CDN, SDN, Q);
   input D, EN, CDN, SDN;
   output Q;
   reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
     buf      (CDN_i, CDN_d);
     buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
     buf      (CDN_i, CDN);
     buf      (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
   not		(E, EN_d);
   tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN_i, notifier);
   buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
   buf      (CDN_i, CDN);
   buf      (SDN_i, SDN);
   not		(E, EN);
   tsmc_dla	(Q_buf, D, E, CDN_i, SDN_i, notifier);
   buf          (Q, Q_buf);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN &&& EN_DEFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
      $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
    $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSNDQD4BWP12TLVT (D, EN, CDN, SDN, Q);
   input D, EN, CDN, SDN;
   output Q;
   reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
     buf      (CDN_i, CDN_d);
     buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
     buf      (CDN_i, CDN);
     buf      (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
   not		(E, EN_d);
   tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN_i, notifier);
   buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
   buf      (CDN_i, CDN);
   buf      (SDN_i, SDN);
   not		(E, EN);
   tsmc_dla	(Q_buf, D, E, CDN_i, SDN_i, notifier);
   buf          (Q, Q_buf);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN &&& EN_DEFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
      $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
    $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSNQD1BWP12TLVT (D, EN, CDN, SDN, Q);
   input D, EN, CDN, SDN;
   output Q;
   reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
     buf      (CDN_i, CDN_d);
     buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
     buf      (CDN_i, CDN);
     buf      (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
   not		(E, EN_d);
   tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN_i, notifier);
   buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
   buf      (CDN_i, CDN);
   buf      (SDN_i, SDN);
   not		(E, EN);
   tsmc_dla	(Q_buf, D, E, CDN_i, SDN_i, notifier);
   buf          (Q, Q_buf);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN &&& EN_DEFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
      $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
    $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSNQD2BWP12TLVT (D, EN, CDN, SDN, Q);
   input D, EN, CDN, SDN;
   output Q;
   reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
     buf      (CDN_i, CDN_d);
     buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
     buf      (CDN_i, CDN);
     buf      (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
   not		(E, EN_d);
   tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN_i, notifier);
   buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
   buf      (CDN_i, CDN);
   buf      (SDN_i, SDN);
   not		(E, EN);
   tsmc_dla	(Q_buf, D, E, CDN_i, SDN_i, notifier);
   buf          (Q, Q_buf);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN &&& EN_DEFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
      $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
    $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSNQD4BWP12TLVT (D, EN, CDN, SDN, Q);
   input D, EN, CDN, SDN;
   output Q;
   reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
     buf      (CDN_i, CDN_d);
     buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
     buf      (CDN_i, CDN);
     buf      (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
   not		(E, EN_d);
   tsmc_dla	(Q_buf, D_d, E, CDN_i, SDN_i, notifier);
   buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
   buf      (CDN_i, CDN);
   buf      (SDN_i, SDN);
   not		(E, EN);
   tsmc_dla	(Q_buf, D, E, CDN_i, SDN_i, notifier);
   buf          (Q, Q_buf);
  `endif
    reg flag;
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  and  (D_check, SDN_i, CDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (CDN => Q) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN, posedge EN &&& EN_DEFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
      $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge CDN, posedge EN &&& EN_DEFCHK, 0, notifier);
    $hold (posedge EN &&& EN_DEFCHK, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LND1BWP12TLVT (D, EN, Q, QN);
    input D, EN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, EN_d ;
    pullup	 (CDN);
    pullup	 (SDN);
    not		 (E, EN_d);
    tsmc_dla (Q_buf, D_d, E, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup	 (CDN);
    pullup	 (SDN);
    not		 (E, EN);
    tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `endif



  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge EN, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge EN, posedge D, 0, 0, notifier,,, EN_d, D_d);
    $setuphold (posedge EN, negedge D, 0, 0, notifier,,, EN_d, D_d);
  `else
    $setuphold (posedge EN, posedge D, 0, 0, notifier);
    $setuphold (posedge EN, negedge D, 0, 0, notifier);
  `endif
  endspecify
endmodule
`endcelldefine

`celldefine
module LND2BWP12TLVT (D, EN, Q, QN);
    input D, EN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, EN_d ;
    pullup	 (CDN);
    pullup	 (SDN);
    not		 (E, EN_d);
    tsmc_dla (Q_buf, D_d, E, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup	 (CDN);
    pullup	 (SDN);
    not		 (E, EN);
    tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `endif



  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge EN, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge EN, posedge D, 0, 0, notifier,,, EN_d, D_d);
    $setuphold (posedge EN, negedge D, 0, 0, notifier,,, EN_d, D_d);
  `else
    $setuphold (posedge EN, posedge D, 0, 0, notifier);
    $setuphold (posedge EN, negedge D, 0, 0, notifier);
  `endif
  endspecify
endmodule
`endcelldefine

`celldefine
module LND4BWP12TLVT (D, EN, Q, QN);
    input D, EN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, EN_d ;
    pullup	 (CDN);
    pullup	 (SDN);
    not		 (E, EN_d);
    tsmc_dla (Q_buf, D_d, E, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup	 (CDN);
    pullup	 (SDN);
    not		 (E, EN);
    tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not		 (QN, Q_buf);
  `endif



  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge EN, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge EN, posedge D, 0, 0, notifier,,, EN_d, D_d);
    $setuphold (posedge EN, negedge D, 0, 0, notifier,,, EN_d, D_d);
  `else
    $setuphold (posedge EN, posedge D, 0, 0, notifier);
    $setuphold (posedge EN, negedge D, 0, 0, notifier);
  `endif
  endspecify
endmodule
`endcelldefine

`celldefine
module LNQD1BWP12TLVT (D, EN, Q);
    input D, EN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, EN_d ;
    pullup	(CDN);
    pullup	(SDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup	(CDN);
    pullup	(SDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge EN, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge EN, posedge D, 0, 0, notifier,,, EN_d, D_d);
    $setuphold (posedge EN, negedge D, 0, 0, notifier,,, EN_d, D_d);
  `else
    $setuphold (posedge EN, posedge D, 0, 0, notifier);
    $setuphold (posedge EN, negedge D, 0, 0, notifier);
  `endif
  endspecify
endmodule
`endcelldefine

`celldefine
module LNQD2BWP12TLVT (D, EN, Q);
    input D, EN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, EN_d ;
    pullup	(CDN);
    pullup	(SDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup	(CDN);
    pullup	(SDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge EN, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge EN, posedge D, 0, 0, notifier,,, EN_d, D_d);
    $setuphold (posedge EN, negedge D, 0, 0, notifier,,, EN_d, D_d);
  `else
    $setuphold (posedge EN, posedge D, 0, 0, notifier);
    $setuphold (posedge EN, negedge D, 0, 0, notifier);
  `endif
  endspecify
endmodule
`endcelldefine

`celldefine
module LNQD4BWP12TLVT (D, EN, Q);
    input D, EN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire D_d, EN_d ;
    pullup	(CDN);
    pullup	(SDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup	(CDN);
    pullup	(SDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge EN, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge EN, posedge D, 0, 0, notifier,,, EN_d, D_d);
    $setuphold (posedge EN, negedge D, 0, 0, notifier,,, EN_d, D_d);
  `else
    $setuphold (posedge EN, posedge D, 0, 0, notifier);
    $setuphold (posedge EN, negedge D, 0, 0, notifier);
  `endif
  endspecify
endmodule
`endcelldefine

`celldefine
module LNSND1BWP12TLVT (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
    pullup       (CDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup       (CDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSND2BWP12TLVT (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
    pullup       (CDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup       (CDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSND4BWP12TLVT (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
    pullup       (CDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup       (CDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSNDD1BWP12TLVT (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
    pullup       (CDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup       (CDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSNDD2BWP12TLVT (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
    pullup       (CDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup       (CDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSNDD4BWP12TLVT (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
    pullup       (CDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup       (CDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
    not		(QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    (SDN => QN) = (0, 0);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSNDQD1BWP12TLVT (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
    pullup       (CDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup       (CDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSNDQD2BWP12TLVT (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
    pullup       (CDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup       (CDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSNDQD4BWP12TLVT (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
    pullup       (CDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup       (CDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSNQD1BWP12TLVT (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
    pullup       (CDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup       (CDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSNQD2BWP12TLVT (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
    pullup       (CDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup       (CDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSNQD4BWP12TLVT (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf          (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (SDN_i, SDN);
    `endif
    wire D_d, EN_d ;
    pullup       (CDN);
    not		(E, EN_d);
    tsmc_dla	(Q_buf, D_d, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (SDN_i, SDN);
    pullup       (CDN);
    not		(E, EN);
    tsmc_dla	(Q_buf, D, E, CDN, SDN_i, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  buf  (D_check, SDN_i);
  buf  (EN_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (SDN => Q) = (0, 0);
    $width (negedge EN, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN, posedge EN, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN, posedge EN, 0, notifier);
      $hold (posedge EN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge EN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $recovery (posedge SDN, posedge EN, 0, notifier);
    $hold (posedge EN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module MAOI222D0BWP12TLVT (A, B, C, ZN);
    input A, B, C;
    output ZN;
    and		(AB, A, B);
    and		(AC, A, C);
    and		(BC, B, C);
    nor		(ZN, AB, AC, BC);

  specify
    (A => ZN) = (0, 0);
    (B => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI222D1BWP12TLVT (A, B, C, ZN);
    input A, B, C;
    output ZN;
    and		(AB, A, B);
    and		(AC, A, C);
    and		(BC, B, C);
    nor		(ZN, AB, AC, BC);

  specify
    (A => ZN) = (0, 0);
    (B => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI222D2BWP12TLVT (A, B, C, ZN);
    input A, B, C;
    output ZN;
    and		(AB, A, B);
    and		(AC, A, C);
    and		(BC, B, C);
    nor		(ZN, AB, AC, BC);

  specify
    (A => ZN) = (0, 0);
    (B => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI222D4BWP12TLVT (A, B, C, ZN);
    input A, B, C;
    output ZN;
    and		(AB, A, B);
    and		(AC, A, C);
    and		(BC, B, C);
    nor		(ZN, AB, AC, BC);

  specify
    (A => ZN) = (0, 0);
    (B => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI22D0BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and		(A, A1, A2);
    nor		(B, B1, B2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI22D1BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and		(A, A1, A2);
    nor		(B, B1, B2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI22D2BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and		(A, A1, A2);
    nor		(B, B1, B2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI22D4BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and		(A, A1, A2);
    nor		(B, B1, B2);
    nor		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MOAI22D0BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or		(A, A1, A2);
    nand		(B, B1, B2);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MOAI22D1BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or		(A, A1, A2);
    nand		(B, B1, B2);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MOAI22D2BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or		(A, A1, A2);
    nand		(B, B1, B2);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MOAI22D4BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or		(A, A1, A2);
    nand		(B, B1, B2);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2D0BWP12TLVT (I0, I1, S, Z);
   input I0, I1, S;
   output Z;
   tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    ifnone (I0 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    ifnone (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
    ifnone (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2D1BWP12TLVT (I0, I1, S, Z);
   input I0, I1, S;
   output Z;
   tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    ifnone (I0 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    ifnone (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
    ifnone (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2D2BWP12TLVT (I0, I1, S, Z);
   input I0, I1, S;
   output Z;
   tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    ifnone (I0 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    ifnone (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
    ifnone (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2D4BWP12TLVT (I0, I1, S, Z);
   input I0, I1, S;
   output Z;
   tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    ifnone (I0 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    ifnone (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
    ifnone (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2ND0BWP12TLVT (I0, I1, S, ZN);
   input I0, I1, S;
   output ZN;
   tsmc_mux (I0_out, I0, I1, S);
   not (ZN, I0_out);

  specify
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    ifnone (I0 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    ifnone (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
    ifnone (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2ND1BWP12TLVT (I0, I1, S, ZN);
   input I0, I1, S;
   output ZN;
   tsmc_mux (I0_out, I0, I1, S);
   not (ZN, I0_out);

  specify
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    ifnone (I0 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    ifnone (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
    ifnone (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2ND2BWP12TLVT (I0, I1, S, ZN);
   input I0, I1, S;
   output ZN;
   tsmc_mux (I0_out, I0, I1, S);
   not (ZN, I0_out);

  specify
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    ifnone (I0 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    ifnone (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
    ifnone (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2ND4BWP12TLVT (I0, I1, S, ZN);
   input I0, I1, S;
   output ZN;
   tsmc_mux (I0_out, I0, I1, S);
   not (ZN, I0_out);

  specify
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    ifnone (I0 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    ifnone (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
    ifnone (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3D0BWP12TLVT (I0, I1, I2, S0, S1, Z);
   input I0, I1, I2, S0, S1;
   output Z;
   tsmc_mux (I0_out, I0, I1, S0);
   tsmc_mux (Z, I0_out, I2, S1);

  specify
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    ifnone (I0 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    ifnone (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    ifnone (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    ifnone (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    ifnone (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3D1BWP12TLVT (I0, I1, I2, S0, S1, Z);
   input I0, I1, I2, S0, S1;
   output Z;
   tsmc_mux (I0_out, I0, I1, S0);
   tsmc_mux (Z, I0_out, I2, S1);

  specify
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    ifnone (I0 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    ifnone (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    ifnone (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    ifnone (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    ifnone (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3D2BWP12TLVT (I0, I1, I2, S0, S1, Z);
   input I0, I1, I2, S0, S1;
   output Z;
   tsmc_mux (I0_out, I0, I1, S0);
   tsmc_mux (Z, I0_out, I2, S1);

  specify
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    ifnone (I0 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    ifnone (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    ifnone (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    ifnone (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    ifnone (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3D4BWP12TLVT (I0, I1, I2, S0, S1, Z);
   input I0, I1, I2, S0, S1;
   output Z;
   tsmc_mux (I0_out, I0, I1, S0);
   tsmc_mux (Z, I0_out, I2, S1);

  specify
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    ifnone (I0 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    ifnone (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    ifnone (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    ifnone (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    ifnone (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3ND0BWP12TLVT (I0, I1, I2, S0, S1, ZN);
   input I0, I1, I2, S0, S1;
   output ZN;
   tsmc_mux (I0_out, I0, I1, S0);
   tsmc_mux (I1_out, I0_out, I2, S1);
   not (ZN, I1_out);

  specify
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    ifnone (I0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    ifnone (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    ifnone (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    ifnone (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    ifnone (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3ND1BWP12TLVT (I0, I1, I2, S0, S1, ZN);
   input I0, I1, I2, S0, S1;
   output ZN;
   tsmc_mux (I0_out, I0, I1, S0);
   tsmc_mux (I1_out, I0_out, I2, S1);
   not (ZN, I1_out);

  specify
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    ifnone (I0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    ifnone (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    ifnone (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    ifnone (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    ifnone (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3ND2BWP12TLVT (I0, I1, I2, S0, S1, ZN);
   input I0, I1, I2, S0, S1;
   output ZN;
   tsmc_mux (I0_out, I0, I1, S0);
   tsmc_mux (I1_out, I0_out, I2, S1);
   not (ZN, I1_out);

  specify
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    ifnone (I0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    ifnone (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    ifnone (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    ifnone (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    ifnone (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3ND4BWP12TLVT (I0, I1, I2, S0, S1, ZN);
   input I0, I1, I2, S0, S1;
   output ZN;
   tsmc_mux (I0_out, I0, I1, S0);
   tsmc_mux (I1_out, I0_out, I2, S1);
   not (ZN, I1_out);

  specify
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    ifnone (I0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    ifnone (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    ifnone (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    ifnone (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    ifnone (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4D0BWP12TLVT (I0, I1, I2, I3, S0, S1, Z);
   input I0, I1, I2, I3, S0, S1;
   output Z;
   tsmc_mux (I0_out, I2, I3, S0);
   tsmc_mux (I1_out, I0, I1, S0);
   tsmc_mux (Z, I1_out, I0_out, S1);

  specify
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    ifnone (I0 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    ifnone (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    ifnone (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    ifnone (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    ifnone (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    ifnone (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4D1BWP12TLVT (I0, I1, I2, I3, S0, S1, Z);
   input I0, I1, I2, I3, S0, S1;
   output Z;
   tsmc_mux (I0_out, I2, I3, S0);
   tsmc_mux (I1_out, I0, I1, S0);
   tsmc_mux (Z, I1_out, I0_out, S1);

  specify
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    ifnone (I0 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    ifnone (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    ifnone (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    ifnone (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    ifnone (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    ifnone (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4D2BWP12TLVT (I0, I1, I2, I3, S0, S1, Z);
   input I0, I1, I2, I3, S0, S1;
   output Z;
   tsmc_mux (I0_out, I2, I3, S0);
   tsmc_mux (I1_out, I0, I1, S0);
   tsmc_mux (Z, I1_out, I0_out, S1);

  specify
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    ifnone (I0 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    ifnone (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    ifnone (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    ifnone (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    ifnone (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    ifnone (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4D4BWP12TLVT (I0, I1, I2, I3, S0, S1, Z);
   input I0, I1, I2, I3, S0, S1;
   output Z;
   tsmc_mux (I0_out, I2, I3, S0);
   tsmc_mux (I1_out, I0, I1, S0);
   tsmc_mux (Z, I1_out, I0_out, S1);

  specify
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    ifnone (I0 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    ifnone (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    ifnone (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    ifnone (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    ifnone (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    ifnone (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4ND0BWP12TLVT (I0, I1, I2, I3, S0, S1, ZN);
   input I0, I1, I2, I3, S0, S1;
   output ZN;
   tsmc_mux (I0_out, I2, I3, S0);
   tsmc_mux (I1_out, I0, I1, S0);
   tsmc_mux (I2_out, I1_out, I0_out, S1);
   not (ZN, I2_out);

  specify
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    ifnone (I0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    ifnone (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    ifnone (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    ifnone (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    ifnone (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    ifnone (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4ND1BWP12TLVT (I0, I1, I2, I3, S0, S1, ZN);
   input I0, I1, I2, I3, S0, S1;
   output ZN;
   tsmc_mux (I0_out, I2, I3, S0);
   tsmc_mux (I1_out, I0, I1, S0);
   tsmc_mux (I2_out, I1_out, I0_out, S1);
   not (ZN, I2_out);

  specify
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    ifnone (I0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    ifnone (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    ifnone (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    ifnone (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    ifnone (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    ifnone (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4ND2BWP12TLVT (I0, I1, I2, I3, S0, S1, ZN);
   input I0, I1, I2, I3, S0, S1;
   output ZN;
   tsmc_mux (I0_out, I2, I3, S0);
   tsmc_mux (I1_out, I0, I1, S0);
   tsmc_mux (I2_out, I1_out, I0_out, S1);
   not (ZN, I2_out);

  specify
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    ifnone (I0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    ifnone (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    ifnone (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    ifnone (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    ifnone (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    ifnone (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4ND4BWP12TLVT (I0, I1, I2, I3, S0, S1, ZN);
   input I0, I1, I2, I3, S0, S1;
   output ZN;
   tsmc_mux (I0_out, I2, I3, S0);
   tsmc_mux (I1_out, I0, I1, S0);
   tsmc_mux (I2_out, I1_out, I0_out, S1);
   not (ZN, I2_out);

  specify
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    ifnone (I0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    ifnone (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    ifnone (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    ifnone (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    ifnone (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    ifnone (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D0BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nand		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D1BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nand		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D2BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nand		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D3BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nand		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D4BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nand		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D8BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nand		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3D0BWP12TLVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    nand		(ZN, A1, A2, A3);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3D1BWP12TLVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    nand		(ZN, A1, A2, A3);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3D2BWP12TLVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    nand		(ZN, A1, A2, A3);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3D3BWP12TLVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    nand		(ZN, A1, A2, A3);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3D4BWP12TLVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    nand		(ZN, A1, A2, A3);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3D8BWP12TLVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    nand		(ZN, A1, A2, A3);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND4D0BWP12TLVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    nand		(ZN, A1, A2, A3, A4);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND4D1BWP12TLVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    nand		(ZN, A1, A2, A3, A4);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND4D2BWP12TLVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    nand		(ZN, A1, A2, A3, A4);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND4D3BWP12TLVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    nand		(ZN, A1, A2, A3, A4);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND4D4BWP12TLVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    nand		(ZN, A1, A2, A3, A4);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND4D8BWP12TLVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    nand		(ZN, A1, A2, A3, A4);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D0BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nor		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D1BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nor		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D2BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nor		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D3BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nor		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D4BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nor		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D8BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nor		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2XD0BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nor		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2XD1BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nor		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2XD2BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nor		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2XD3BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nor		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2XD4BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nor		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2XD8BWP12TLVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    nor		(ZN, A1, A2);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3D0BWP12TLVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    nor		(ZN, A1, A2, A3);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3D1BWP12TLVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    nor		(ZN, A1, A2, A3);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3D2BWP12TLVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    nor		(ZN, A1, A2, A3);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3D3BWP12TLVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    nor		(ZN, A1, A2, A3);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3D4BWP12TLVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    nor		(ZN, A1, A2, A3);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3D8BWP12TLVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    nor		(ZN, A1, A2, A3);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR4D0BWP12TLVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    nor		(ZN, A1, A2, A3, A4);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR4D1BWP12TLVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    nor		(ZN, A1, A2, A3, A4);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR4D2BWP12TLVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    nor		(ZN, A1, A2, A3, A4);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR4D3BWP12TLVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    nor		(ZN, A1, A2, A3, A4);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR4D4BWP12TLVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    nor		(ZN, A1, A2, A3, A4);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR4D8BWP12TLVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    nor		(ZN, A1, A2, A3, A4);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA211D0BWP12TLVT (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    or		(A, A1, A2);
    and		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B => Z) = (0, 0);
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA211D1BWP12TLVT (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    or		(A, A1, A2);
    and		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B => Z) = (0, 0);
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA211D2BWP12TLVT (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    or		(A, A1, A2);
    and		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B => Z) = (0, 0);
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA211D4BWP12TLVT (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    or		(A, A1, A2);
    and		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B => Z) = (0, 0);
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA21D0BWP12TLVT (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    or		(A, A1, A2);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA21D1BWP12TLVT (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    or		(A, A1, A2);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA21D2BWP12TLVT (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    or		(A, A1, A2);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA21D4BWP12TLVT (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    or		(A, A1, A2);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA221D0BWP12TLVT (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    or		(A, A1, A2);
    or      (B, B1, B2);
    and		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA221D1BWP12TLVT (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    or		(A, A1, A2);
    or      (B, B1, B2);
    and		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA221D2BWP12TLVT (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    or		(A, A1, A2);
    or      (B, B1, B2);
    and		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA221D4BWP12TLVT (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    or		(A, A1, A2);
    or      (B, B1, B2);
    and		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA222D0BWP12TLVT (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    or		(A, A1, A2);
    or      (B, B1, B2);
    or      (C, C1, C2);
    and		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (C1 => Z) = (0, 0);
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA222D1BWP12TLVT (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    or		(A, A1, A2);
    or      (B, B1, B2);
    or      (C, C1, C2);
    and		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (C1 => Z) = (0, 0);
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA222D2BWP12TLVT (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    or		(A, A1, A2);
    or      (B, B1, B2);
    or      (C, C1, C2);
    and		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (C1 => Z) = (0, 0);
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA222D4BWP12TLVT (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    or		(A, A1, A2);
    or      (B, B1, B2);
    or      (C, C1, C2);
    and		(Z, A, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (C1 => Z) = (0, 0);
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA22D0BWP12TLVT (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    or		(A, A1, A2);
    or      (B, B1, B2);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA22D1BWP12TLVT (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    or		(A, A1, A2);
    or      (B, B1, B2);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA22D2BWP12TLVT (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    or		(A, A1, A2);
    or      (B, B1, B2);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA22D4BWP12TLVT (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    or		(A, A1, A2);
    or      (B, B1, B2);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA31D0BWP12TLVT (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    or		(A, A1, A2, A3);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA31D1BWP12TLVT (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    or		(A, A1, A2, A3);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA31D2BWP12TLVT (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    or		(A, A1, A2, A3);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA31D4BWP12TLVT (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    or		(A, A1, A2, A3);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA32D0BWP12TLVT (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    or		(A, A1, A2, A3);
    or		(B, B1, B2);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA32D1BWP12TLVT (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    or		(A, A1, A2, A3);
    or		(B, B1, B2);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA32D2BWP12TLVT (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    or		(A, A1, A2, A3);
    or		(B, B1, B2);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA32D4BWP12TLVT (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    or		(A, A1, A2, A3);
    or		(B, B1, B2);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA33D0BWP12TLVT (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    or		(A, A1, A2, A3);
    or		(B, B1, B2, B3);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA33D1BWP12TLVT (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    or		(A, A1, A2, A3);
    or		(B, B1, B2, B3);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA33D2BWP12TLVT (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    or		(A, A1, A2, A3);
    or		(B, B1, B2, B3);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA33D4BWP12TLVT (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    or		(A, A1, A2, A3);
    or		(B, B1, B2, B3);
    and		(Z, A, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (B1 => Z) = (0, 0);
    (B2 => Z) = (0, 0);
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI211D0BWP12TLVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    or		(A, A1, A2);
    nand		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI211D1BWP12TLVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    or		(A, A1, A2);
    nand		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI211D2BWP12TLVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    or		(A, A1, A2);
    nand		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI211D4BWP12TLVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    or		(A, A1, A2);
    nand		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI21D0BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or		(A, A1, A2);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI21D1BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or		(A, A1, A2);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI21D2BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or		(A, A1, A2);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI21D4BWP12TLVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or		(A, A1, A2);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI221D0BWP12TLVT (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    or		(A, A1, A2);
    or		(B, B1, B2);
    nand         (ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI221D1BWP12TLVT (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    or		(A, A1, A2);
    or		(B, B1, B2);
    nand         (ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI221D2BWP12TLVT (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    or		(A, A1, A2);
    or		(B, B1, B2);
    nand         (ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI221D4BWP12TLVT (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    or		(A, A1, A2);
    or		(B, B1, B2);
    nand         (ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI221XD4BWP12TLVT (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    or		(A, A1, A2);
    or		(B, B1, B2);
    nand         (ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI222D0BWP12TLVT (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    or		(A, A1, A2);
    or		(B, B1, B2);
    or		(C, C1, C2);
    nand		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C1 => ZN) = (0, 0);
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI222D1BWP12TLVT (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    or		(A, A1, A2);
    or		(B, B1, B2);
    or		(C, C1, C2);
    nand		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C1 => ZN) = (0, 0);
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI222D2BWP12TLVT (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    or		(A, A1, A2);
    or		(B, B1, B2);
    or		(C, C1, C2);
    nand		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C1 => ZN) = (0, 0);
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI222D4BWP12TLVT (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    or		(A, A1, A2);
    or		(B, B1, B2);
    or		(C, C1, C2);
    nand		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C1 => ZN) = (0, 0);
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI222XD4BWP12TLVT (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    or		(A, A1, A2);
    or		(B, B1, B2);
    or		(C, C1, C2);
    nand		(ZN, A, B, C);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (C1 => ZN) = (0, 0);
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI22D0BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or		(A, A1, A2);
    or		(B, B1, B2);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI22D1BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or		(A, A1, A2);
    or		(B, B1, B2);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI22D2BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or		(A, A1, A2);
    or		(B, B1, B2);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI22D4BWP12TLVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or		(A, A1, A2);
    or		(B, B1, B2);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI31D0BWP12TLVT (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    or		(A, A1, A2, A3);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI31D1BWP12TLVT (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    or		(A, A1, A2, A3);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI31D2BWP12TLVT (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    or		(A, A1, A2, A3);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI31D4BWP12TLVT (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    or		(A, A1, A2, A3);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI32D0BWP12TLVT (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    or		(A, A1, A2, A3);
    or		(B, B1, B2);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI32D1BWP12TLVT (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    or		(A, A1, A2, A3);
    or		(B, B1, B2);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI32D2BWP12TLVT (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    or		(A, A1, A2, A3);
    or		(B, B1, B2);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI32D4BWP12TLVT (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    or		(A, A1, A2, A3);
    or		(B, B1, B2);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI32XD4BWP12TLVT (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    or		(A, A1, A2, A3);
    or		(B, B1, B2);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI33D0BWP12TLVT (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    or		(A, A1, A2, A3);
    or		(B, B1, B2, B3);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI33D1BWP12TLVT (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    or		(A, A1, A2, A3);
    or		(B, B1, B2, B3);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI33D2BWP12TLVT (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    or		(A, A1, A2, A3);
    or		(B, B1, B2, B3);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI33D4BWP12TLVT (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    or		(A, A1, A2, A3);
    or		(B, B1, B2, B3);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI33XD4BWP12TLVT (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    or		(A, A1, A2, A3);
    or		(B, B1, B2, B3);
    nand		(ZN, A, B);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OD25DCAP16BWP12TLVT;
    // No function
endmodule
`endcelldefine

`celldefine
module OD25DCAP32BWP12TLVT;
    // No function
endmodule
`endcelldefine

`celldefine
module OD25DCAP64BWP12TLVT;
    // No function
endmodule
`endcelldefine

`celldefine
module OR2D0BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2D1BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2D2BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2D4BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2D8BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2XD1BWP12TLVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or		(Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR3D0BWP12TLVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    or		(Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR3D1BWP12TLVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    or		(Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR3D2BWP12TLVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    or		(Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR3D4BWP12TLVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    or		(Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR3D8BWP12TLVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    or		(Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR3XD1BWP12TLVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    or		(Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR4D0BWP12TLVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    or		(Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR4D1BWP12TLVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    or		(Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR4D2BWP12TLVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    or		(Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR4D4BWP12TLVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    or		(Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR4D8BWP12TLVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    or		(Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR4XD1BWP12TLVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    or		(Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module SDFCND0BWP12TLVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    pullup   (SDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    pullup   (SDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CP_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCND1BWP12TLVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    pullup   (SDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    pullup   (SDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CP_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCND2BWP12TLVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    pullup   (SDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    pullup   (SDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CP_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCND4BWP12TLVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    pullup   (SDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    pullup   (SDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CP_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNQD0BWP12TLVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    pullup       (SDN);
    tsmc_mux     (D_i, D_d, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CP_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNQD1BWP12TLVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    pullup       (SDN);
    tsmc_mux     (D_i, D_d, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CP_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNQD2BWP12TLVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    pullup       (SDN);
    tsmc_mux     (D_i, D_d, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CP_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNQD4BWP12TLVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf          (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf          (CDN_i, CDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    pullup       (SDN);
    tsmc_mux     (D_i, D_d, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf          (CDN_i, CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN_i, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CP_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSND0BWP12TLVT (SI, D, SE, CP, CDN, SDN, Q, QN);
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    reg flag;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `endif
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CP_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSND1BWP12TLVT (SI, D, SE, CP, CDN, SDN, Q, QN);
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    reg flag;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `endif
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CP_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSND2BWP12TLVT (SI, D, SE, CP, CDN, SDN, Q, QN);
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    reg flag;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `endif
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CP_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSND4BWP12TLVT (SI, D, SE, CP, CDN, SDN, Q, QN);
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    reg flag;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `endif
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CP_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSNQD0BWP12TLVT (SI, D, SE, CP, CDN, SDN, Q);
    input SI, D, SE, CP, CDN, SDN;
    output Q;
    reg notifier;
    reg flag;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CP_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSNQD1BWP12TLVT (SI, D, SE, CP, CDN, SDN, Q);
    input SI, D, SE, CP, CDN, SDN;
    output Q;
    reg notifier;
    reg flag;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CP_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSNQD2BWP12TLVT (SI, D, SE, CP, CDN, SDN, Q);
    input SI, D, SE, CP, CDN, SDN;
    output Q;
    reg notifier;
    reg flag;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CP_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSNQD4BWP12TLVT (SI, D, SE, CP, CDN, SDN, Q);
    input SI, D, SE, CP, CDN, SDN;
    output Q;
    reg notifier;
    reg flag;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CP_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFD0BWP12TLVT (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D_d, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFD1BWP12TLVT (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D_d, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFD2BWP12TLVT (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D_d, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFD4BWP12TLVT (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D_d, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCND0BWP12TLVT (SI, D, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d ;
    pullup   (CDN);
    pullup   (SDN);
    and      (D1, CN_d, D_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    and      (D1, CN, D);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCND1BWP12TLVT (SI, D, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d ;
    pullup   (CDN);
    pullup   (SDN);
    and      (D1, CN_d, D_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    and      (D1, CN, D);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCND2BWP12TLVT (SI, D, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d ;
    pullup   (CDN);
    pullup   (SDN);
    and      (D1, CN_d, D_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    and      (D1, CN, D);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCND4BWP12TLVT (SI, D, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d ;
    pullup   (CDN);
    pullup   (SDN);
    and      (D1, CN_d, D_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    and      (D1, CN, D);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCNQD0BWP12TLVT (SI, D, SE, CP, CN, Q);
    input SI, D, SE, CP, CN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d ;
    pullup (CDN);
    pullup (SDN);
    and (D1, CN_d, D_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup (CDN);
    pullup (SDN);
    and (D1, CN, D);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCNQD1BWP12TLVT (SI, D, SE, CP, CN, Q);
    input SI, D, SE, CP, CN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d ;
    pullup (CDN);
    pullup (SDN);
    and (D1, CN_d, D_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup (CDN);
    pullup (SDN);
    and (D1, CN, D);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCNQD2BWP12TLVT (SI, D, SE, CP, CN, Q);
    input SI, D, SE, CP, CN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d ;
    pullup (CDN);
    pullup (SDN);
    and (D1, CN_d, D_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup (CDN);
    pullup (SDN);
    and (D1, CN, D);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCNQD4BWP12TLVT (SI, D, SE, CP, CN, Q);
    input SI, D, SE, CP, CN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d ;
    pullup (CDN);
    pullup (SDN);
    and (D1, CN_d, D_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup (CDN);
    pullup (SDN);
    and (D1, CN, D);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSND0BWP12TLVT (SI, D, SE, CP, CN, SN, Q, QN);
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d ;
    pullup (CDN); 
    pullup (SDN);
    not (S, SN_d);
    or  (DS, S, D_d);
    and (D1, DS, CN_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);  
    buf (Q, Q_buf);        
    not (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup (CDN); 
    pullup (SDN);
    not (S, SN);
    or  (DS, S, D);
    and (D1, DS, CN);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);  
    buf (Q, Q_buf);        
    not (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d, SN_d);
    and  (SN_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN, SN);
    and  (SN_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSND1BWP12TLVT (SI, D, SE, CP, CN, SN, Q, QN);
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d ;
    pullup (CDN); 
    pullup (SDN);
    not (S, SN_d);
    or  (DS, S, D_d);
    and (D1, DS, CN_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);  
    buf (Q, Q_buf);        
    not (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup (CDN); 
    pullup (SDN);
    not (S, SN);
    or  (DS, S, D);
    and (D1, DS, CN);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);  
    buf (Q, Q_buf);        
    not (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d, SN_d);
    and  (SN_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN, SN);
    and  (SN_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSND2BWP12TLVT (SI, D, SE, CP, CN, SN, Q, QN);
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d ;
    pullup (CDN); 
    pullup (SDN);
    not (S, SN_d);
    or  (DS, S, D_d);
    and (D1, DS, CN_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);  
    buf (Q, Q_buf);        
    not (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup (CDN); 
    pullup (SDN);
    not (S, SN);
    or  (DS, S, D);
    and (D1, DS, CN);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);  
    buf (Q, Q_buf);        
    not (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d, SN_d);
    and  (SN_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN, SN);
    and  (SN_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSND4BWP12TLVT (SI, D, SE, CP, CN, SN, Q, QN);
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d ;
    pullup (CDN); 
    pullup (SDN);
    not (S, SN_d);
    or  (DS, S, D_d);
    and (D1, DS, CN_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);  
    buf (Q, Q_buf);        
    not (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup (CDN); 
    pullup (SDN);
    not (S, SN);
    or  (DS, S, D);
    and (D1, DS, CN);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);  
    buf (Q, Q_buf);        
    not (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d, SN_d);
    and  (SN_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN, SN);
    and  (SN_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSNQD0BWP12TLVT (SI, D, SE, CP, CN, SN, Q);
    input SI, D, SE, CP, CN, SN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d ;
    pullup (CDN); 
    pullup (SDN);
    not (S, SN_d);
    or  (DS, S, D_d);
    and (D1, DS, CN_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);  
    buf (Q, Q_buf);        
  `else 	// Reserve for non NTC.
    pullup (CDN); 
    pullup (SDN);
    not (S, SN);
    or  (DS, S, D);
    and (D1, DS, CN);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);  
    buf (Q, Q_buf);        
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d, SN_d);
    and  (SN_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN, SN);
    and  (SN_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSNQD1BWP12TLVT (SI, D, SE, CP, CN, SN, Q);
    input SI, D, SE, CP, CN, SN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d ;
    pullup (CDN); 
    pullup (SDN);
    not (S, SN_d);
    or  (DS, S, D_d);
    and (D1, DS, CN_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);  
    buf (Q, Q_buf);        
  `else 	// Reserve for non NTC.
    pullup (CDN); 
    pullup (SDN);
    not (S, SN);
    or  (DS, S, D);
    and (D1, DS, CN);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);  
    buf (Q, Q_buf);        
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d, SN_d);
    and  (SN_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN, SN);
    and  (SN_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSNQD2BWP12TLVT (SI, D, SE, CP, CN, SN, Q);
    input SI, D, SE, CP, CN, SN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d ;
    pullup (CDN); 
    pullup (SDN);
    not (S, SN_d);
    or  (DS, S, D_d);
    and (D1, DS, CN_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);  
    buf (Q, Q_buf);        
  `else 	// Reserve for non NTC.
    pullup (CDN); 
    pullup (SDN);
    not (S, SN);
    or  (DS, S, D);
    and (D1, DS, CN);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);  
    buf (Q, Q_buf);        
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d, SN_d);
    and  (SN_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN, SN);
    and  (SN_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSNQD4BWP12TLVT (SI, D, SE, CP, CN, SN, Q);
    input SI, D, SE, CP, CN, SN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d ;
    pullup (CDN); 
    pullup (SDN);
    not (S, SN_d);
    or  (DS, S, D_d);
    and (D1, DS, CN_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);  
    buf (Q, Q_buf);        
  `else 	// Reserve for non NTC.
    pullup (CDN); 
    pullup (SDN);
    not (S, SN);
    or  (DS, S, D);
    and (D1, DS, CN);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);  
    buf (Q, Q_buf);        
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, CN_d, SN_d);
    and  (SN_check, SE_int_not, CN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, CN, SN);
    and  (SN_check, SE_int_not, CN);
  `endif
  buf  (CN_check, SE_int_not);
   `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSND0BWP12TLVT (SI, D, SE, CP, SN, Q, QN);
    input SI, D, SE, CP, SN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, SN_d ;
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN_d);     
    or       (D1, S, D_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN);     
    or       (D1, S, D);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, SN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, SN);
  `endif
  buf  (SN_check, SE_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSND1BWP12TLVT (SI, D, SE, CP, SN, Q, QN);
    input SI, D, SE, CP, SN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, SN_d ;
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN_d);     
    or       (D1, S, D_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN);     
    or       (D1, S, D);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, SN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, SN);
  `endif
  buf  (SN_check, SE_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSND2BWP12TLVT (SI, D, SE, CP, SN, Q, QN);
    input SI, D, SE, CP, SN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, SN_d ;
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN_d);     
    or       (D1, S, D_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN);     
    or       (D1, S, D);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, SN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, SN);
  `endif
  buf  (SN_check, SE_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSND4BWP12TLVT (SI, D, SE, CP, SN, Q, QN);
    input SI, D, SE, CP, SN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, SN_d ;
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN_d);     
    or       (D1, S, D_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN);     
    or       (D1, S, D);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, SN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, SN);
  `endif
  buf  (SN_check, SE_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSNQD0BWP12TLVT (SI, D, SE, CP, SN, Q);
    input SI, D, SE, CP, SN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, SN_d ;
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN_d);     
    or       (D1, S, D_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
  `else 	// Reserve for non NTC.
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN);     
    or       (D1, S, D);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, SN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, SN);
  `endif
  buf  (SN_check, SE_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSNQD1BWP12TLVT (SI, D, SE, CP, SN, Q);
    input SI, D, SE, CP, SN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, SN_d ;
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN_d);     
    or       (D1, S, D_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
  `else 	// Reserve for non NTC.
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN);     
    or       (D1, S, D);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, SN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, SN);
  `endif
  buf  (SN_check, SE_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSNQD2BWP12TLVT (SI, D, SE, CP, SN, Q);
    input SI, D, SE, CP, SN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, SN_d ;
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN_d);     
    or       (D1, S, D_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
  `else 	// Reserve for non NTC.
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN);     
    or       (D1, S, D);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, SN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, SN);
  `endif
  buf  (SN_check, SE_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSNQD4BWP12TLVT (SI, D, SE, CP, SN, Q);
    input SI, D, SE, CP, SN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, SN_d ;
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN_d);     
    or       (D1, S, D_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
  `else 	// Reserve for non NTC.
    pullup   (CDN); 
    pullup   (SDN);
    not      (S, SN);     
    or       (D1, S, D);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);  
    buf      (Q, Q_buf);        
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, SE_int_not, SN_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, SE_int_not, SN);
  `endif
  buf  (SN_check, SE_int_not);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP, 0, 0, notifier);
    $width (negedge CP, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, posedge SN, 0, 0, notifier);
    $setuphold (posedge CP &&& SN_DEFCHK, negedge SN, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCND0BWP12TLVT (SI, D, SE, CPN, CDN, Q, QN);
    input SI, D, SE, CPN, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire SI_d, D_d, SE_d, CPN_d ;
    pullup   (SDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    not      (CP, CPN_d);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    pullup   (SDN);
    tsmc_mux (D_i, D, SI, SE);
    not      (CP, CPN);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CPN_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN, negedge CPN, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCND1BWP12TLVT (SI, D, SE, CPN, CDN, Q, QN);
    input SI, D, SE, CPN, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire SI_d, D_d, SE_d, CPN_d ;
    pullup   (SDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    not      (CP, CPN_d);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    pullup   (SDN);
    tsmc_mux (D_i, D, SI, SE);
    not      (CP, CPN);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CPN_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN, negedge CPN, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCND2BWP12TLVT (SI, D, SE, CPN, CDN, Q, QN);
    input SI, D, SE, CPN, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire SI_d, D_d, SE_d, CPN_d ;
    pullup   (SDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    not      (CP, CPN_d);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    pullup   (SDN);
    tsmc_mux (D_i, D, SI, SE);
    not      (CP, CPN);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CPN_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN, negedge CPN, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCND4BWP12TLVT (SI, D, SE, CPN, CDN, Q, QN);
    input SI, D, SE, CPN, CDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire SI_d, D_d, SE_d, CPN_d ;
    pullup   (SDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    not      (CP, CPN_d);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    pullup   (SDN);
    tsmc_mux (D_i, D, SI, SE);
    not      (CP, CPN);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
  `endif
  and  (D_check, CDN_i, SE_int_not);
  buf  (CPN_check, CDN_i);
  buf  (SE_check, CDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN, negedge CPN, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCSND0BWP12TLVT (SI, D, SE, CPN, CDN, SDN, Q, QN);
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    reg flag;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CPN_d ;
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    not	     (CP, CPN_d);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_mux (D_i, D, SI, SE);
    not	     (CP, CPN);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `endif
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CPN_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN, negedge CPN, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, negedge CPN, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCSND1BWP12TLVT (SI, D, SE, CPN, CDN, SDN, Q, QN);
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    reg flag;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CPN_d ;
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    not	     (CP, CPN_d);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_mux (D_i, D, SI, SE);
    not	     (CP, CPN);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `endif
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CPN_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN, negedge CPN, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, negedge CPN, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCSND2BWP12TLVT (SI, D, SE, CPN, CDN, SDN, Q, QN);
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    reg flag;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CPN_d ;
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    not	     (CP, CPN_d);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_mux (D_i, D, SI, SE);
    not	     (CP, CPN);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `endif
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CPN_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN, negedge CPN, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, negedge CPN, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCSND4BWP12TLVT (SI, D, SE, CPN, CDN, SDN, Q, QN);
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    reg flag;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d , SDN_d ;
      buf      (CDN_i, CDN_d);
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CPN_d ;
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    not	     (CP, CPN_d);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `else 	// Reserve for non NTC.
    buf      (CDN_i, CDN);
    buf      (SDN_i, SDN);
    tsmc_mux (D_i, D, SI, SE);
    not	     (CP, CPN);
    tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN_buf, Q_buf);
    and      (QN, QN_buf, SDN_i);
  `endif
    always @(CDN_i or SDN_i) begin
      if (!$test$plusargs("cdn_sdn_check_off")) begin
      if (flag == 1) begin 
         if (CDN_i!==1'b0) begin
         $display("%m > CDN is released at time %.2fns.", $realtime);
         end
         if (SDN_i!==1'b0) begin
         $display("%m > SDN is released at time %.2fns.", $realtime);
         end
      end
      flag = ((CDN_i===1'b0)&&(SDN_i ===1'b0));
      if (flag == 1) begin
         $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
      end
    end 
    end



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SDN_i, SE);
  `endif
  and  (D_check, CDN_i, SDN_i, SE_int_not);
  and  (CPN_check, CDN_i, SDN_i);
  and  (SE_check, CDN_i, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN, negedge CPN, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN, posedge SDN, 0,0, notifier, , , CDN_d, SDN_d);
      $recrem (posedge SDN, negedge CPN, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN, posedge CDN, 0,0, notifier, , , SDN_d, CDN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge CDN, 0, notifier);
      $recovery (posedge CDN, posedge SDN, 0, notifier);
      $hold (posedge SDN, posedge CDN, 0, notifier);
      $recovery (posedge SDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge SDN, 0, notifier);
      $recovery (posedge SDN, posedge CDN, 0, notifier);
      $hold (posedge CDN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge CDN, 0, notifier);
    $recovery (posedge CDN, posedge SDN, 0, notifier);
    $hold (posedge SDN, posedge CDN, 0, notifier);
    $recovery (posedge SDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge SDN, 0, notifier);
    $recovery (posedge SDN, posedge CDN, 0, notifier);
    $hold (posedge CDN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFND0BWP12TLVT (SI, D, SE, CPN, Q, QN);
    input SI, D, SE, CPN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CPN_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D_d, SI_d, SE_d);
    not		 (CP, CPN_d);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D, SI, SE);
    not		 (CP, CPN);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CPN_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFND1BWP12TLVT (SI, D, SE, CPN, Q, QN);
    input SI, D, SE, CPN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CPN_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D_d, SI_d, SE_d);
    not		 (CP, CPN_d);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D, SI, SE);
    not		 (CP, CPN);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CPN_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFND2BWP12TLVT (SI, D, SE, CPN, Q, QN);
    input SI, D, SE, CPN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CPN_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D_d, SI_d, SE_d);
    not		 (CP, CPN_d);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D, SI, SE);
    not		 (CP, CPN);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CPN_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFND4BWP12TLVT (SI, D, SE, CPN, Q, QN);
    input SI, D, SE, CPN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CPN_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D_d, SI_d, SE_d);
    not		 (CP, CPN_d);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D, SI, SE);
    not		 (CP, CPN);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CPN_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSND0BWP12TLVT (SI, D, SE, CPN, SDN, Q, QN);
    input SI, D, SE, CPN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CPN_d ;
    pullup   (CDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    not	     (CP, CPN_d);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (SDN_i, SDN);
    pullup   (CDN);
    tsmc_mux (D_i, D, SI, SE);
    not	     (CP, CPN);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CPN_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge SDN, negedge CPN, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge SDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge SDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSND1BWP12TLVT (SI, D, SE, CPN, SDN, Q, QN);
    input SI, D, SE, CPN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CPN_d ;
    pullup   (CDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    not	     (CP, CPN_d);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (SDN_i, SDN);
    pullup   (CDN);
    tsmc_mux (D_i, D, SI, SE);
    not	     (CP, CPN);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CPN_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge SDN, negedge CPN, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge SDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge SDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSND2BWP12TLVT (SI, D, SE, CPN, SDN, Q, QN);
    input SI, D, SE, CPN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CPN_d ;
    pullup   (CDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    not	     (CP, CPN_d);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (SDN_i, SDN);
    pullup   (CDN);
    tsmc_mux (D_i, D, SI, SE);
    not	     (CP, CPN);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CPN_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge SDN, negedge CPN, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge SDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge SDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSND4BWP12TLVT (SI, D, SE, CPN, SDN, Q, QN);
    input SI, D, SE, CPN, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CPN_d ;
    pullup   (CDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    not	     (CP, CPN_d);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (SDN_i, SDN);
    pullup   (CDN);
    tsmc_mux (D_i, D, SI, SE);
    not	     (CP, CPN);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CPN_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CPN_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge SDN, negedge CPN, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge SDN, negedge CPN, 0, notifier);
      $hold (negedge CPN, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (negedge CPN &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge SDN, negedge CPN, 0, notifier);
    $hold (negedge CPN, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQD0BWP12TLVT (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQD1BWP12TLVT (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQD2BWP12TLVT (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQD4BWP12TLVT (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQND0BWP12TLVT (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D_d, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    not          (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    not          (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQND1BWP12TLVT (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D_d, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    not          (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    not          (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQND2BWP12TLVT (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D_d, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    not          (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    not          (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQND4BWP12TLVT (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D_d, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    not          (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    not          (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
  `else
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
  `endif
  buf  (D_check, SE_int_not);
  pullup  (CP_check);
  pullup  (SE_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSND0BWP12TLVT (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    pullup   (CDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (SDN_i, SDN);
    pullup   (CDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CP_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSND1BWP12TLVT (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    pullup   (CDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (SDN_i, SDN);
    pullup   (CDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CP_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSND2BWP12TLVT (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    pullup   (CDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (SDN_i, SDN);
    pullup   (CDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CP_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSND4BWP12TLVT (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    pullup   (CDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (SDN_i, SDN);
    pullup   (CDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CP_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSNQD0BWP12TLVT (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    pullup   (CDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (SDN_i, SDN);
    pullup   (CDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CP_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSNQD1BWP12TLVT (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    pullup   (CDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (SDN_i, SDN);
    pullup   (CDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CP_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSNQD2BWP12TLVT (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    pullup   (CDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (SDN_i, SDN);
    pullup   (CDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CP_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSNQD4BWP12TLVT (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  SDN_d ;
      buf      (SDN_i, SDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (SDN_i, SDN);
    `endif
    wire SI_d, D_d, SE_d, CP_d ;
    pullup   (CDN);
    tsmc_mux (D_i, D_d, SI_d, SE_d);
    tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    buf      (SDN_i, SDN);
    pullup   (CDN);
    tsmc_mux (D_i, D, SI, SE);
    tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SE_int_not, SE_d);
    and  (SI_check, SDN_i, SE_d);
  `else
    not  (SE_int_not, SE);
    and  (SI_check, SDN_i, SE);
  `endif
  and  (D_check, SDN_i, SE_int_not);
  buf  (CP_check, SDN_i);
  buf  (SE_check, SDN_i);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge SDN, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN, posedge CP, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge SDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SE_DEFCHK, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge SDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge SDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFXD0BWP12TLVT (DA, DB, SA, SI, SE, CP, Q, QN);
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB_d, DA_d, SA_d);
    tsmc_mux     (D_i, D, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB, DA, SA);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (DA_check, SA_d, SE_int_not);
  `else
    not  (SA_int_not, SA);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (DA_check, SA, SE_int_not);
  `endif
  buf  (SA_check, SE_int_not);
  and  (DB_check, SA_int_not, SE_int_not);
  or   (CP_check, SI_check, DA_check, SA_check, DB_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFXD1BWP12TLVT (DA, DB, SA, SI, SE, CP, Q, QN);
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB_d, DA_d, SA_d);
    tsmc_mux     (D_i, D, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB, DA, SA);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (DA_check, SA_d, SE_int_not);
  `else
    not  (SA_int_not, SA);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (DA_check, SA, SE_int_not);
  `endif
  buf  (SA_check, SE_int_not);
  and  (DB_check, SA_int_not, SE_int_not);
  or   (CP_check, SI_check, DA_check, SA_check, DB_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFXD2BWP12TLVT (DA, DB, SA, SI, SE, CP, Q, QN);
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB_d, DA_d, SA_d);
    tsmc_mux     (D_i, D, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB, DA, SA);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (DA_check, SA_d, SE_int_not);
  `else
    not  (SA_int_not, SA);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (DA_check, SA, SE_int_not);
  `endif
  buf  (SA_check, SE_int_not);
  and  (DB_check, SA_int_not, SE_int_not);
  or   (CP_check, SI_check, DA_check, SA_check, DB_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFXD4BWP12TLVT (DA, DB, SA, SI, SE, CP, Q, QN);
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB_d, DA_d, SA_d);
    tsmc_mux     (D_i, D, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB, DA, SA);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
    not          (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (DA_check, SA_d, SE_int_not);
  `else
    not  (SA_int_not, SA);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (DA_check, SA, SE_int_not);
  `endif
  buf  (SA_check, SE_int_not);
  and  (DB_check, SA_int_not, SE_int_not);
  or   (CP_check, SI_check, DA_check, SA_check, DB_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFXQD0BWP12TLVT (DA, DB, SA, SI, SE, CP, Q);
    input DA, DB, SA, SI, SE, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB_d, DA_d, SA_d);
    tsmc_mux     (D_i, D, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB, DA, SA);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (DA_check, SA_d, SE_int_not);
  `else
    not  (SA_int_not, SA);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (DA_check, SA, SE_int_not);
  `endif
  buf  (SA_check, SE_int_not);
  and  (DB_check, SA_int_not, SE_int_not);
  or   (CP_check, SI_check, DA_check, SA_check, DB_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFXQD1BWP12TLVT (DA, DB, SA, SI, SE, CP, Q);
    input DA, DB, SA, SI, SE, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB_d, DA_d, SA_d);
    tsmc_mux     (D_i, D, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB, DA, SA);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (DA_check, SA_d, SE_int_not);
  `else
    not  (SA_int_not, SA);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (DA_check, SA, SE_int_not);
  `endif
  buf  (SA_check, SE_int_not);
  and  (DB_check, SA_int_not, SE_int_not);
  or   (CP_check, SI_check, DA_check, SA_check, DB_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFXQD2BWP12TLVT (DA, DB, SA, SI, SE, CP, Q);
    input DA, DB, SA, SI, SE, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB_d, DA_d, SA_d);
    tsmc_mux     (D_i, D, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB, DA, SA);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (DA_check, SA_d, SE_int_not);
  `else
    not  (SA_int_not, SA);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (DA_check, SA, SE_int_not);
  `endif
  buf  (SA_check, SE_int_not);
  and  (DB_check, SA_int_not, SE_int_not);
  or   (CP_check, SI_check, DA_check, SA_check, DB_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFXQD4BWP12TLVT (DA, DB, SA, SI, SE, CP, Q);
    input DA, DB, SA, SI, SE, CP;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d ;
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB_d, DA_d, SA_d);
    tsmc_mux     (D_i, D, SI_d, SE_d);
    tsmc_dff     (Q_buf, D_i, CP_d, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup       (CDN);
    pullup       (SDN);
    tsmc_mux     (D, DB, DA, SA);
    tsmc_mux     (D_i, D, SI, SE);
    tsmc_dff     (Q_buf, D_i, CP, CDN, SDN, notifier);
    buf          (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (SA_int_not, SA_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (DA_check, SA_d, SE_int_not);
  `else
    not  (SA_int_not, SA);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (DA_check, SA, SE_int_not);
  `endif
  buf  (SA_check, SE_int_not);
  and  (DB_check, SA_int_not, SE_int_not);
  or   (CP_check, SI_check, DA_check, SA_check, DB_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DA_DEFCHK, posedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DEFCHK, negedge DA, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, posedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& DB_DEFCHK, negedge DB, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, posedge SA, 0, 0, notifier);
    $setuphold (posedge CP &&& SA_DEFCHK, negedge SA, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFCND0BWP12TLVT (E, SE, CP, SI, D, CDN, Q, QN);
    input E, SE, CP, SI, D, CDN; 
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (SDN);
    buf      (CDN_i, CDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
    and  (D_check, CDN_i, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
    and  (D_check, CDN_i, E, SE_int_not);
  `endif
  and  (E_check, CDN_i, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFCND1BWP12TLVT (E, SE, CP, SI, D, CDN, Q, QN);
    input E, SE, CP, SI, D, CDN; 
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (SDN);
    buf      (CDN_i, CDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
    and  (D_check, CDN_i, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
    and  (D_check, CDN_i, E, SE_int_not);
  `endif
  and  (E_check, CDN_i, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFCND2BWP12TLVT (E, SE, CP, SI, D, CDN, Q, QN);
    input E, SE, CP, SI, D, CDN; 
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (SDN);
    buf      (CDN_i, CDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
    and  (D_check, CDN_i, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
    and  (D_check, CDN_i, E, SE_int_not);
  `endif
  and  (E_check, CDN_i, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFCND4BWP12TLVT (E, SE, CP, SI, D, CDN, Q, QN);
    input E, SE, CP, SI, D, CDN; 
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (SDN);
    buf      (CDN_i, CDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
    and  (D_check, CDN_i, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
    and  (D_check, CDN_i, E, SE_int_not);
  `endif
  and  (E_check, CDN_i, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFCNQD0BWP12TLVT (E, SE, CP, SI, D, CDN, Q);
    input E, SE, CP, SI, D, CDN; 
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (SDN);
    buf      (CDN_i, CDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
    and  (D_check, CDN_i, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
    and  (D_check, CDN_i, E, SE_int_not);
  `endif
  and  (E_check, CDN_i, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFCNQD1BWP12TLVT (E, SE, CP, SI, D, CDN, Q);
    input E, SE, CP, SI, D, CDN; 
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (SDN);
    buf      (CDN_i, CDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
    and  (D_check, CDN_i, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
    and  (D_check, CDN_i, E, SE_int_not);
  `endif
  and  (E_check, CDN_i, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFCNQD2BWP12TLVT (E, SE, CP, SI, D, CDN, Q);
    input E, SE, CP, SI, D, CDN; 
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (SDN);
    buf      (CDN_i, CDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
    and  (D_check, CDN_i, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
    and  (D_check, CDN_i, E, SE_int_not);
  `endif
  and  (E_check, CDN_i, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFCNQD4BWP12TLVT (E, SE, CP, SI, D, CDN, Q);
    input E, SE, CP, SI, D, CDN; 
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    `ifdef RECREM 	// Reserve for RECREM.
      wire  CDN_d ;
      buf      (CDN_i, CDN_d);
    `else         	// Reserve for non RECREM. 
      buf      (CDN_i, CDN);
    `endif
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (SDN);
    buf      (CDN_i, CDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN_i, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (SI_check, CDN_i, SE_d);
    and  (D_check, CDN_i, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (SI_check, CDN_i, SE);
    and  (D_check, CDN_i, E, SE_int_not);
  `endif
  and  (E_check, CDN_i, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (negedge CDN, 0, 0, notifier);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN, posedge CP, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
      $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN, posedge CP, 0, notifier);
      $hold (posedge CP, posedge CDN, 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
    $recovery (posedge CDN, posedge CP, 0, notifier);
    $hold (posedge CP, posedge CDN, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFD0BWP12TLVT (E, SE, CP, SI, D, Q, QN);
    input E, SE, CP, SI, D; 
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFD1BWP12TLVT (E, SE, CP, SI, D, Q, QN);
    input E, SE, CP, SI, D; 
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFD2BWP12TLVT (E, SE, CP, SI, D, Q, QN);
    input E, SE, CP, SI, D; 
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFD4BWP12TLVT (E, SE, CP, SI, D, Q, QN);
    input E, SE, CP, SI, D; 
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFKCND0BWP12TLVT (SI, D, E, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN, E;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d, E_d ;
    pullup (CDN);
    pullup (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    and (D2, CN_d, D1);
    tsmc_mux (D3, D2, SI_d, SE_d);
    tsmc_dff (Q_buf, D3, CP_d, CDN, SDN, notifier);
    buf (Q, Q_buf);
    not (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup (CDN);
    pullup (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    and (D2, CN, D1);
    tsmc_mux (D3, D2, SI, SE);
    tsmc_dff (Q_buf, D3, CP, CDN, SDN, notifier);
    buf (Q, Q_buf);
    not (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (D_check, E_d, CN_d, SE_int_not);
    and  (E_check, CN_d, SE_int_not);
    buf  (SI_check, SE_d);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (D_check, E, CN, SE_int_not);
    and  (E_check, CN, SE_int_not);
    buf  (SI_check, SE);
  `endif
  buf  (CN_check, SE_int_not);
  or   (CP_check, D_check, E_check, CN_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFKCND1BWP12TLVT (SI, D, E, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN, E;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d, E_d ;
    pullup (CDN);
    pullup (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    and (D2, CN_d, D1);
    tsmc_mux (D3, D2, SI_d, SE_d);
    tsmc_dff (Q_buf, D3, CP_d, CDN, SDN, notifier);
    buf (Q, Q_buf);
    not (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup (CDN);
    pullup (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    and (D2, CN, D1);
    tsmc_mux (D3, D2, SI, SE);
    tsmc_dff (Q_buf, D3, CP, CDN, SDN, notifier);
    buf (Q, Q_buf);
    not (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (D_check, E_d, CN_d, SE_int_not);
    and  (E_check, CN_d, SE_int_not);
    buf  (SI_check, SE_d);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (D_check, E, CN, SE_int_not);
    and  (E_check, CN, SE_int_not);
    buf  (SI_check, SE);
  `endif
  buf  (CN_check, SE_int_not);
  or   (CP_check, D_check, E_check, CN_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFKCND2BWP12TLVT (SI, D, E, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN, E;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d, E_d ;
    pullup (CDN);
    pullup (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    and (D2, CN_d, D1);
    tsmc_mux (D3, D2, SI_d, SE_d);
    tsmc_dff (Q_buf, D3, CP_d, CDN, SDN, notifier);
    buf (Q, Q_buf);
    not (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup (CDN);
    pullup (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    and (D2, CN, D1);
    tsmc_mux (D3, D2, SI, SE);
    tsmc_dff (Q_buf, D3, CP, CDN, SDN, notifier);
    buf (Q, Q_buf);
    not (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (D_check, E_d, CN_d, SE_int_not);
    and  (E_check, CN_d, SE_int_not);
    buf  (SI_check, SE_d);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (D_check, E, CN, SE_int_not);
    and  (E_check, CN, SE_int_not);
    buf  (SI_check, SE);
  `endif
  buf  (CN_check, SE_int_not);
  or   (CP_check, D_check, E_check, CN_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFKCND4BWP12TLVT (SI, D, E, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN, E;
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d, E_d ;
    pullup (CDN);
    pullup (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    and (D2, CN_d, D1);
    tsmc_mux (D3, D2, SI_d, SE_d);
    tsmc_dff (Q_buf, D3, CP_d, CDN, SDN, notifier);
    buf (Q, Q_buf);
    not (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup (CDN);
    pullup (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    and (D2, CN, D1);
    tsmc_mux (D3, D2, SI, SE);
    tsmc_dff (Q_buf, D3, CP, CDN, SDN, notifier);
    buf (Q, Q_buf);
    not (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (D_check, E_d, CN_d, SE_int_not);
    and  (E_check, CN_d, SE_int_not);
    buf  (SI_check, SE_d);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (D_check, E, CN, SE_int_not);
    and  (E_check, CN, SE_int_not);
    buf  (SI_check, SE);
  `endif
  buf  (CN_check, SE_int_not);
  or   (CP_check, D_check, E_check, CN_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFKCNQD0BWP12TLVT (SI, D, E, SE, CP, CN, Q);
    input SI, D, SE, CP, CN, E;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d, E_d ;
    pullup (CDN);
    pullup (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    and (D2, CN_d, D1);
    tsmc_mux (D3, D2, SI_d, SE_d);
    tsmc_dff (Q_buf, D3, CP_d, CDN, SDN, notifier);
    buf (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup (CDN);
    pullup (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    and (D2, CN, D1);
    tsmc_mux (D3, D2, SI, SE);
    tsmc_dff (Q_buf, D3, CP, CDN, SDN, notifier);
    buf (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (D_check, E_d, CN_d, SE_int_not);
    and  (E_check, CN_d, SE_int_not);
    buf  (SI_check, SE_d);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (D_check, E, CN, SE_int_not);
    and  (E_check, CN, SE_int_not);
    buf  (SI_check, SE);
  `endif
  buf  (CN_check, SE_int_not);
  or   (CP_check, D_check, E_check, CN_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFKCNQD1BWP12TLVT (SI, D, E, SE, CP, CN, Q);
    input SI, D, SE, CP, CN, E;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d, E_d ;
    pullup (CDN);
    pullup (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    and (D2, CN_d, D1);
    tsmc_mux (D3, D2, SI_d, SE_d);
    tsmc_dff (Q_buf, D3, CP_d, CDN, SDN, notifier);
    buf (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup (CDN);
    pullup (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    and (D2, CN, D1);
    tsmc_mux (D3, D2, SI, SE);
    tsmc_dff (Q_buf, D3, CP, CDN, SDN, notifier);
    buf (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (D_check, E_d, CN_d, SE_int_not);
    and  (E_check, CN_d, SE_int_not);
    buf  (SI_check, SE_d);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (D_check, E, CN, SE_int_not);
    and  (E_check, CN, SE_int_not);
    buf  (SI_check, SE);
  `endif
  buf  (CN_check, SE_int_not);
  or   (CP_check, D_check, E_check, CN_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFKCNQD2BWP12TLVT (SI, D, E, SE, CP, CN, Q);
    input SI, D, SE, CP, CN, E;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d, E_d ;
    pullup (CDN);
    pullup (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    and (D2, CN_d, D1);
    tsmc_mux (D3, D2, SI_d, SE_d);
    tsmc_dff (Q_buf, D3, CP_d, CDN, SDN, notifier);
    buf (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup (CDN);
    pullup (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    and (D2, CN, D1);
    tsmc_mux (D3, D2, SI, SE);
    tsmc_dff (Q_buf, D3, CP, CDN, SDN, notifier);
    buf (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (D_check, E_d, CN_d, SE_int_not);
    and  (E_check, CN_d, SE_int_not);
    buf  (SI_check, SE_d);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (D_check, E, CN, SE_int_not);
    and  (E_check, CN, SE_int_not);
    buf  (SI_check, SE);
  `endif
  buf  (CN_check, SE_int_not);
  or   (CP_check, D_check, E_check, CN_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFKCNQD4BWP12TLVT (SI, D, E, SE, CP, CN, Q);
    input SI, D, SE, CP, CN, E;
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire SI_d, D_d, SE_d, CP_d, CN_d, E_d ;
    pullup (CDN);
    pullup (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    and (D2, CN_d, D1);
    tsmc_mux (D3, D2, SI_d, SE_d);
    tsmc_dff (Q_buf, D3, CP_d, CDN, SDN, notifier);
    buf (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup (CDN);
    pullup (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    and (D2, CN, D1);
    tsmc_mux (D3, D2, SI, SE);
    tsmc_dff (Q_buf, D3, CP, CDN, SDN, notifier);
    buf (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    and  (D_check, E_d, CN_d, SE_int_not);
    and  (E_check, CN_d, SE_int_not);
    buf  (SI_check, SE_d);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    and  (D_check, E, CN, SE_int_not);
    and  (E_check, CN, SE_int_not);
    buf  (SI_check, SE);
  `endif
  buf  (CN_check, SE_int_not);
  or   (CP_check, D_check, E_check, CN_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && E && D) || (!(SE) && CN && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& CN_DEFCHK, posedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& CN_DEFCHK, negedge CN, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQD0BWP12TLVT (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D; 
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQD1BWP12TLVT (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D; 
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQD2BWP12TLVT (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D; 
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQD4BWP12TLVT (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D; 
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQND0BWP12TLVT (E, SE, CP, SI, D, QN);
    input E, SE, CP, SI, D; 
    output QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQND1BWP12TLVT (E, SE, CP, SI, D, QN);
    input E, SE, CP, SI, D; 
    output QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQND2BWP12TLVT (E, SE, CP, SI, D, QN);
    input E, SE, CP, SI, D; 
    output QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQND4BWP12TLVT (E, SE, CP, SI, D, QN);
    input E, SE, CP, SI, D; 
    output QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQNXD0BWP12TLVT (E, SE, CP, SI, D, QN);
    input E, SE, CP, SI, D; 
    output QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQNXD1BWP12TLVT (E, SE, CP, SI, D, QN);
    input E, SE, CP, SI, D; 
    output QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQNXD2BWP12TLVT (E, SE, CP, SI, D, QN);
    input E, SE, CP, SI, D; 
    output QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQNXD4BWP12TLVT (E, SE, CP, SI, D, QN);
    input E, SE, CP, SI, D; 
    output QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQXD0BWP12TLVT (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D; 
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQXD1BWP12TLVT (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D; 
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQXD2BWP12TLVT (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D; 
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFQXD4BWP12TLVT (E, SE, CP, SI, D, Q);
    input E, SE, CP, SI, D; 
    output Q;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFXD0BWP12TLVT (E, SE, CP, SI, D, Q, QN);
    input E, SE, CP, SI, D; 
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFXD1BWP12TLVT (E, SE, CP, SI, D, Q, QN);
    input E, SE, CP, SI, D; 
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFXD2BWP12TLVT (E, SE, CP, SI, D, Q, QN);
    input E, SE, CP, SI, D; 
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SEDFXD4BWP12TLVT (E, SE, CP, SI, D, Q, QN);
    input E, SE, CP, SI, D; 
    output Q, QN;
    reg notifier;
  `ifdef NTC 	// Reserve for NTC.
    wire E_d, SE_d, CP_d, SI_d, D_d ;
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D_d, E_d);
    tsmc_mux (D2, D1, SI_d, SE_d);
    tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `else 	// Reserve for non NTC.
    pullup   (CDN);
    pullup   (SDN);
    tsmc_mux (D1, Q_buf, D, E);
    tsmc_mux (D2, D1, SI, SE);
    tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
    buf      (Q, Q_buf);
    not      (QN, Q_buf);
  `endif



  // Timing logics defined for default constraint check
  `ifdef NTC
    not  (E_int_not, E_d);
    not  (SE_int_not, SE_d);
    buf  (SI_check, SE_d);
    and  (D_check, E_d, SE_int_not);
  `else
    not  (E_int_not, E);
    not  (SE_int_not, SE);
    buf  (SI_check, SE);
    and  (D_check, E, SE_int_not);
  `endif
  buf  (E_check, SE_int_not);
  or   (CP_check, D_check, E_check, SI_check);
  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
  `endif

  `ifdef TETRAMAX
  `else
  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && E && D) || (!(SE) && !(E) && Q_buf)))) = (0, 0);
    $width (posedge CP &&& CP_DEFCHK, 0, 0, notifier);
    $width (negedge CP &&& CP_DEFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, posedge E, 0, 0, notifier);
    $setuphold (posedge CP &&& E_DEFCHK, negedge E, 0, 0, notifier);
    $setuphold (posedge CP, posedge SE, 0, 0, notifier);
    $setuphold (posedge CP, negedge SE, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, posedge SI, 0, 0, notifier);
    $setuphold (posedge CP &&& SI_DEFCHK, negedge SI, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module TIEHBWP12TLVT (Z);
  output  Z;
  buf (Z, 1'b1);

endmodule
`endcelldefine

`celldefine
module TIELBWP12TLVT (ZN);
  output  ZN;
  buf (ZN, 1'b0);

endmodule
`endcelldefine

`celldefine
module XNR2D0BWP12TLVT (A1, A2, ZN);
  input		A1, A2;
  output 	ZN;
  xnor		(ZN, A1, A2);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    ifnone (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
    ifnone (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR2D1BWP12TLVT (A1, A2, ZN);
  input		A1, A2;
  output 	ZN;
  xnor		(ZN, A1, A2);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    ifnone (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
    ifnone (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR2D2BWP12TLVT (A1, A2, ZN);
  input		A1, A2;
  output 	ZN;
  xnor		(ZN, A1, A2);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    ifnone (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
    ifnone (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR2D4BWP12TLVT (A1, A2, ZN);
  input		A1, A2;
  output 	ZN;
  xnor		(ZN, A1, A2);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    ifnone (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
    ifnone (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR3D0BWP12TLVT (A1, A2, A3, ZN);
  input A1, A2, A3;
  output ZN;
  xnor		(ZN, A1, A2, A3);

  specify
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    ifnone (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    ifnone (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    ifnone (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR3D1BWP12TLVT (A1, A2, A3, ZN);
  input A1, A2, A3;
  output ZN;
  xnor		(ZN, A1, A2, A3);

  specify
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    ifnone (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    ifnone (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    ifnone (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR3D2BWP12TLVT (A1, A2, A3, ZN);
  input A1, A2, A3;
  output ZN;
  xnor		(ZN, A1, A2, A3);

  specify
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    ifnone (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    ifnone (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    ifnone (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR3D4BWP12TLVT (A1, A2, A3, ZN);
  input A1, A2, A3;
  output ZN;
  xnor		(ZN, A1, A2, A3);

  specify
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    ifnone (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    ifnone (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    ifnone (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR4D0BWP12TLVT (A1, A2, A3, A4, ZN);
  input 	A1, A2, A3, A4;
  output 	ZN;
  xnor		(ZN, A1, A2, A3, A4);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    ifnone (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    ifnone (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    ifnone (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    ifnone (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR4D1BWP12TLVT (A1, A2, A3, A4, ZN);
  input 	A1, A2, A3, A4;
  output 	ZN;
  xnor		(ZN, A1, A2, A3, A4);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    ifnone (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    ifnone (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    ifnone (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    ifnone (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR4D2BWP12TLVT (A1, A2, A3, A4, ZN);
  input 	A1, A2, A3, A4;
  output 	ZN;
  xnor		(ZN, A1, A2, A3, A4);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    ifnone (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    ifnone (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    ifnone (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    ifnone (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR4D4BWP12TLVT (A1, A2, A3, A4, ZN);
  input 	A1, A2, A3, A4;
  output 	ZN;
  xnor		(ZN, A1, A2, A3, A4);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    ifnone (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    ifnone (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    ifnone (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    ifnone (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR2D0BWP12TLVT (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
  xor		(Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    ifnone (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
    ifnone (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR2D1BWP12TLVT (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
  xor		(Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    ifnone (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
    ifnone (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR2D2BWP12TLVT (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
  xor		(Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    ifnone (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
    ifnone (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR2D4BWP12TLVT (A1, A2, Z);
  input 	A1, A2;
  output 	Z;
  xor		(Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    ifnone (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
    ifnone (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR3D0BWP12TLVT (A1, A2, A3, Z);
  input A1, A2, A3;
  output Z;
  xor		(Z, A1, A2, A3);

  specify
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    ifnone (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    ifnone (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    ifnone (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR3D1BWP12TLVT (A1, A2, A3, Z);
  input A1, A2, A3;
  output Z;
  xor		(Z, A1, A2, A3);

  specify
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    ifnone (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    ifnone (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    ifnone (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR3D2BWP12TLVT (A1, A2, A3, Z);
  input A1, A2, A3;
  output Z;
  xor		(Z, A1, A2, A3);

  specify
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    ifnone (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    ifnone (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    ifnone (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR3D4BWP12TLVT (A1, A2, A3, Z);
  input A1, A2, A3;
  output Z;
  xor		(Z, A1, A2, A3);

  specify
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    ifnone (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    ifnone (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    ifnone (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR4D0BWP12TLVT (A1, A2, A3, A4, Z);
  input 	A1, A2, A3, A4;
  output 	Z;
  xor		(Z, A1, A2, A3, A4);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    ifnone (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    ifnone (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    ifnone (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    ifnone (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR4D1BWP12TLVT (A1, A2, A3, A4, Z);
  input 	A1, A2, A3, A4;
  output 	Z;
  xor		(Z, A1, A2, A3, A4);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    ifnone (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    ifnone (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    ifnone (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    ifnone (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR4D2BWP12TLVT (A1, A2, A3, A4, Z);
  input 	A1, A2, A3, A4;
  output 	Z;
  xor		(Z, A1, A2, A3, A4);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    ifnone (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    ifnone (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    ifnone (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    ifnone (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR4D4BWP12TLVT (A1, A2, A3, A4, Z);
  input 	A1, A2, A3, A4;
  output 	Z;
  xor		(Z, A1, A2, A3, A4);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    ifnone (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    ifnone (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    ifnone (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    ifnone (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOHID1BWP12TLVT (ISO, I, Z);
    input ISO, I;
    output Z;
    or		(Z,I,ISO);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOHID2BWP12TLVT (ISO, I, Z);
    input ISO, I;
    output Z;
    or          (Z,I,ISO);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOHID4BWP12TLVT (ISO, I, Z);
    input ISO, I;
    output Z;
    or          (Z,I,ISO);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOHID8BWP12TLVT (ISO, I, Z);
    input ISO, I;
    output Z;
    or          (Z,I,ISO);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOLOD1BWP12TLVT (ISO, I, Z);
    input ISO, I;
    output Z;
    not		(ISO1, ISO);
    nand	(Z1, ISO1, I);
    not		(Z, Z1);    

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOLOD2BWP12TLVT (ISO, I, Z);
    input ISO, I;
    output Z;
    not         (ISO1, ISO);
    nand        (Z1, ISO1, I);
    not         (Z, Z1);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOLOD4BWP12TLVT (ISO, I, Z);
    input ISO, I;
    output Z;
    not         (ISO1, ISO);
    nand        (Z1, ISO1, I);
    not         (Z, Z1);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOLOD8BWP12TLVT (ISO, I, Z);
    input ISO, I;
    output Z;
    not         (ISO1, ISO);
    nand        (Z1, ISO1, I);
    not         (Z, Z1);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLHLD1BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLHLD2BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLHLD4BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLHLD8BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHCD1BWP12TLVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    not		(IN, I);
    nand		(Z, IN, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHCD2BWP12TLVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    not		(IN, I);
    nand		(Z, IN, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHCD4BWP12TLVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    not		(IN, I);
    nand		(Z, IN, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHCD8BWP12TLVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    not		(IN, I);
    nand		(Z, IN, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHD1BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHD2BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHD4BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHD8BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHFACD1BWP12TLVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    not		(IN, I);
    nand		(Z, IN, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHFACD2BWP12TLVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    not		(IN, I);
    nand		(Z, IN, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHFACD4BWP12TLVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    not		(IN, I);
    nand		(Z, IN, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHFACD8BWP12TLVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    not		(IN, I);
    nand		(Z, IN, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHFACLOD1BWP12TLVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    and		(Z, I, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHFACLOD2BWP12TLVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    and		(Z, I, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHFACLOD4BWP12TLVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    and		(Z, I, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHFACLOD8BWP12TLVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    and		(Z, I, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHFAD1BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHFAD2BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHFAD4BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHFAD8BWP12TLVT (I, Z);
    input I;
    output Z;
    buf		(Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine





primitive tsmc_mux (q, d0, d1, s);
   output q;
   input s, d0, d1;

   table
   // d0  d1  s   : q 
      0   ?   0   : 0 ;
      1   ?   0   : 1 ;
      ?   0   1   : 0 ;
      ?   1   1   : 1 ;
      0   0   x   : 0 ;
      1   1   x   : 1 ;
   endtable
endprimitive
primitive tsmc_dla (q, d, e, cdn, sdn, notifier);
   output q;
   reg q;
   input d, e, cdn, sdn, notifier;
   table
   1  1   1   ?   ?   : ?  :  1  ; // Latch 1
   0  1   ?   1   ?   : ?  :  0  ; // Latch 0
   0 (10) 1   1   ?   : ?  :  0  ; // Latch 0 after falling edge
   1 (10) 1   1   ?   : ?  :  1  ; // Latch 1 after falling edge
   *  0   ?   ?   ?   : ?  :  -  ; // no changes
   ?  ?   ?   0   ?   : ?  :  1  ; // preset to 1
   ?  0   1   *   ?   : 1  :  1  ;
   1  ?   1   *   ?   : 1  :  1  ;
   1  *   1   ?   ?   : 1  :  1  ;
   ?  ?   0   1   ?   : ?  :  0  ; // reset to 0
   ?  0   *   1   ?   : 0  :  0  ;
   0  ?   *   1   ?   : 0  :  0  ;
   0  *   ?   1   ?   : 0  :  0  ;
   ?  ?   ?   ?   *   : ?  :  x  ; // toggle notifier
   endtable
endprimitive
primitive tsmc_xbuf (o, i, dummy);
   output o;     
   input i, dummy;
   table         
   // i dummy : o
      0   1   : 0 ;
      1   1   : 1 ;
      x   1   : 1 ;
   endtable      
endprimitive 
primitive tsmc_dff (q, d, cp, cdn, sdn, notifier);
   output q;
   input d, cp, cdn, sdn, notifier;
   reg q;
   table
      ?   ?   0   ?   ? : ? : 0 ; // CDN dominate SDN
      ?   ?   1   0   ? : ? : 1 ; // SDN is set   
      ?   ?   1   x   ? : 0 : x ; // SDN affect Q
      ?   ?   1   x   ? : 1 : 1 ; // Q=1,preset=X
      ?   ?   x   1   ? : 0 : 0 ; // Q=0,clear=X
      0 (01)  ?   1   ? : ? : 0 ; // Latch 0
      0   *   ?   1   ? : 0 : 0 ; // Keep 0 (D==Q)
      1 (01)  1   ?   ? : ? : 1 ; // Latch 1   
      1   *   1   ?   ? : 1 : 1 ; // Keep 1 (D==Q)
      ? (1?)  1   1   ? : ? : - ; // ignore negative edge of clock
      ? (?0)  1   1   ? : ? : - ; // ignore negative edge of clock
      ?   ? (?1)  1   ? : ? : - ; // ignore positive edge of CDN
      ?   ?   1 (?1)  ? : ? : - ; // ignore posative edge of SDN
      *   ?   1   1   ? : ? : - ; // ignore data change on steady clock
      ?   ?   ?   ?   * : ? : x ; // timing check violation
   endtable
endprimitive
